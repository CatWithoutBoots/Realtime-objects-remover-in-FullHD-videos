��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&r�F���oh���[ynnf���6_�h�0�Kh�G� ��>�.�������4�i��u�ɞ��P���W_�&ML�چ�-�G^Ew$7�����d+9�,��r�"1�*�OلG0��A�<���E�3��Wˆ��V��C�8�0�
���>��m8C��s��!��wZ��
�C���ؼ�Moؙ'�����S�j��p��q�*9��a'�5%'ϥTj���|갃ϸ2�nE���R��W��_��;d���l�0�������[[%H�d��t�c�
{���C.���o����IH`�.at��q�Ѡ�(w��o&@���M��EIZP�
q�EҶ��*˦�5V���I�J�!�Ы��'p-rB����Pyf�#N��iF�.��f:6}���ZئQ�����\BXlP<ةy�$�M���JGe����܁����w�v�����'��޺�Ē�����
$�S?;5`�2$:cn����d�
)�k�t^�4���򎮢���Rp,hM�%:K�k�q�2�p`X0S9��<V�C΋�s���sҘ�Z��$է&�k�N�#�Q�w*P:���wn�ʲ����q��򙻎�}���hi��牏�Ho�2~�u�&$m���c������'�0%�}�m���)�FM���r�y�]�=�]�\�?������˖4��^��I��b�q1��]aT��k<����.VyU#OMr+m7����)Aټ�D�AŴ�_�(�h�r|�ϫ�4��eA�b�o�z�ΐU�'�[k��ǟ�Up��.����Ιݲ�������Y:��k�kD�|@��cr���O��3�����ϩ���Sù "���ۻ��+�_J�\��v���("*a�g��J��;��g���/�[��(���
��(�Q�#m��F���q��fYӦ)��m�� /�'84EΧ4'��E�>��ܴ�['z�dB���}5A_���ѝm)�r���0��VSוs̒�q�zV�ure�UQ+��4���m�'�"��Ŀ|=�J��.�TM��h���HF�!�6��߃�Ũ_��F�e*�.O���o�M�mX��3�+N�'�����b=��<�t��7k�A�Љ�U��p'j����5
�y���"]�ȗZT�W'��O9r<g�87ұ��f.Ei��a D|����[��'r��{_�=�6%�����b�;� �s����19UW�������k&X�����.	ު��Wې�~b�c�g1�w�t+��G����Ŀ���'��q^�n��]���@s�Pv�h�;\�ŋ2��@�उBT1�Z��}VxCl�Ň��E����L-X&w����\��!�~JJt��|������w�=&b�&*��E!�ce�l�)ݥJn/*� t�;��lo�F�D��֤#�k-+���'[����]��t���������a����	�O���S�<B)�ͳ�����ֳf�L��_sꛠyB՜��\�$����q� �b�~�FD섍��2�m�-ˍ����:��Z����T~�����$"V+:QoQp���7ʊﲓ�m�6��	��Tx�x���mZ��Daj@�8(��Q֫���:n	�gW���ı��M���l���{�O�	�|P����焐��u����	3��d��0hK�.��ֻǨ.7u�>���s��j��sN�����	P�X���)	�AC�]W�4#a���V�BT�=%*Y�Gdr�VE6�����.N��Y�Y�������٬�P����X�(�b�� <x�Ǩ��`�4ѓ��?�b �s�������&Wm)_��=|p����'+e��C"0����S��е�{'�:b��6�_���(��ht��b�6��U�b��x����}-[�GG���$�5����hl��ʙS�l�a�(�xzKˋTY��Dj-�@��a���U�K����d�o�{���#��rnk"�!Ew��Hq���R�L�l�N��~:� t�v�Y�m'(�bx9�2}��צ޵T;&�K[��9k���G2����d���_�W�������:�"t�"��@��sU�_1���c�*���K2����y�۟�9z�
�e�� �2(����<�:yw ��J�Pxl/��w�9T��'9��h@�@Q`HčPP:%�o�g�W|�c���UWu���7�����`&6�k?œMğ�Q��Q�4'�Ex:Cb����=�8[�b�po��g?��%{�@����#�Dlq1�Mk��ږ�p�߼iR��=F������U8r�U`.U���(Ԟ�Z�2�S��U�3�n	�F���y�^|�٭��*rt��!b\�ymS�nH�;���B�=�2��!')|��{Mg�y����Q�P �U+�w��cO�,���H��}�B���{O��.;���Bu��`���^u/��m&���vj7&m�M��g�
����gm�GyDʞE�k񏢌uXg����������ؖkS�an�k(gJr���p�$Tm�4(U�Y���Bvs�<���l�c˃)���'Mm�=��;�
�x�d���:�]�%�"�׷���=���f�4sk�"�7W��1c��������|��A�Q�ac�HK�.rm
���q1�ߊ�q�x&d�|y�njuI�3$3�W�0��f��d!���q��孝GI�=��t3�p�eao�#���pρ]O�21^�zaf<�'�H=t5�'������X��7��� �.6>��K]g����O�@�Ӫr����N��<r��;�G{��h�B=���51x�+uwѣ�Y�:H�;!�0k=O���G�i�6��
'GsR�ڡ��֌��x�5��.7��)'�E�@h���˸ #���j���b���0N~ ����=Oe�Kd~@�����\�ze��!��w�L��Tp��\u�\.�:��$�@����+[$�w{w�E5����q��	�r�����-�-_(��:Y Zo��4���66+�݊��A[s��n�Uu�zUO�_C��`QH���9+~���V\v��
�|�ʫr��z��y��Y�SM�%���tv=��&J��I�3f�Vݳ�iS�j[���䑢g,�9��Ў�Xo~�6c�
nx���ƈ��`B[):ĳK���W9V?�"�[��f���MM�R	�d�m���V����2\�C6�`CmQ���2�(<����C��ѥɹ�g �1�!wP�`|^��a�v�o�lj0�\�5*zcڻ��n+����Ux��a�z��#C8ۺR��4�8���� ���\}��n	��4S}ʾ	��݋����֟�������HJ7��ض;4�������g���4��_ԶZ�Z4x���6�����rd�nLݱ����㾗�~��"�O|G�_������y��X�ݻ^�w��O����aF�3嗮�I�H���P���U�ɧ�ou5h���h��pU �iN`��U$P�B?�i�&(.b�%�Z��r4�����s�"�K��~��s���ׁr��0���u���Z�p������Z~��H����=��zd'�!�ؔ�&o,^���Y+��=4�o� ����X*�4�p�H�]��e�u��ѴuO��O/D�����<.����b�8���F'�*���r{�P}Y")�
�U2��9��X@9`��I�{�FP�d��ZC׈��˙T�賞:�@3�0_Ѓ �?8��FN��޻W�X��`78�$(]s:���@�h�ԍ.!eTХŰ��}Ԥ���B�"[�i��2��5�P����Ԭ��<�氅5n$���:����ٙ|����!��p��G^�v��m�b5�M7��h���,m,{\�$@�'R; �F�I*�c���F<&oˣ���N�"y��-U[�!ه�5�h�}�l����L7�$<�����a��abDҽ2uXvT�R[�>������� ���$�b'���|���+�b4'��X	�
�~�+i>��g�x��ԥ���� ���<�8�ne�b��QA$�ƭU��� ���3�;�{���ޤ�i�����au���x�`�7A9�}�C��Y-)��zʅ��"��Ɠ�"f��i�K�+p�'XՋ����p��S�hZ�8��/f63pHo����۵��֌�mKj��g2R�Iu��mʪ)���� 8z��\�ƪ��/�(��|��K^�C��&�z5��@�ܷQr��]�J9�hwT05n��U�;��hY�mT�l�){��p�015����/��,�[&2K�.�)e�� M��C���7���ޭ��Z:ݤFh|�_�Ɵ
�n��r�t�E	���Ҍ_��p�T!�&T|9�1ג�5�h��Z�����j��w�@����2��m���M�c��$�rI�J�q��-)0c��i�ݠH	�X/����}�+�n���hp��@*�f��iDĵ���r�X��e-s�Y��B ��_���F+w`%c�̀��z�Վ�u� �r���f
ۼz�p��P�Bz!�tQeB+���b(�?0ݳ�~�6�_5z�����6	�ZM:cr��~@�g�ӽ�OoȈW�|(��g�6��fa,��		l���I�T�C 
�2�I�\�������s�JB��PS�G���,��o6�p�	�,���f]k��C�ٓ��Z(�v�ܐG�`T�u�� �Yàq��9!�ZVF����i����iL>,<�wI/�w"���G�lJ��j��H��~%��55&l�E�i�ޝ޺o9)2Tޗ�Uez�c:�~>�<6�V�Ƴ���M~��h������iy�#��%L�.j���@�#*�+�%SJ��{f��K�q���E�_r����ضM��wJ�B�W��q/p>�n���&Xko-(L��ZH8'z?T>��T���x���<A�`;ZpQy�@z�9wM���h�D�avhyp*��1�y�0�o�QS
�O�;|�XV;�%?�צ(�TF�A�prc�%�S:nb"��ī����r5�Y��Pҭ������%�M���ﱾ����i����Nfk.��_���Nw��X̥�T���9l�2���ZAbA�^?Ζ6� 2U��g���B��2��I��&�ήm���N.n��1�t���Px�������L�cԷB��UA�- ������ o�j�0�����������/e�xS���$B��h��T�i�"�+���`�"[(o;<O$�glAL�wb���A�9P?EZ`TY�8�&N6}|&��;�[�ھ���`P��8
�ۨ<��2�k�d�~�kկ��_�N�j�U	<w��J<ģ9\Z Z�ZA�aNx��g�f>�뉓���"�Kk���*������r��Vx�"����5�)�}�UĮΞ�6� ��٬�UU�w\)M��H�P����9�s�#�*�|����/Le��[k�t�g����$��� �������o��7;#݋jSS~vJ v� a�����)|b��"
�k{��ŕo�Lz�z�%6�3�F��	�秹 ����f` �
�W�ئ���G��Cw7���v��� ����Z'��5Y��z�-u�`ƫl� Pa�pY��fI��#�������<�w�����%O}�8`0p�I�A����gz^qY�a������LN��|'�N���ן�͇��Ȑۤª�w�L�f�����������rB�-H�1wl�wA%X��Jm��"7^r���n����6?�,��'��b���M� �Z�3��9�Ћ������D���~GĨg�]��#�rJ�X/&a�V0��^� ��)�ʻG�g����j���L^�����B�@ܢ��珐�Dk��Q>L��)����Q�������m X���������i(WGQ�L�mNN�M�0�D��	r�j�ԸZ�f�5���4���/=�C�178���P^~7�o�x"�"Q���K����lA�`T:'���f}�hy�&�2,3��&}�y����e��;e;��w��WW�>�l{{e0���5s���)�u#z�rC9Yߡ;�aUS�A��._K��
J

*.X{�a�ؚ�')~������DMf�f�Ŗ�F��;�1��y�k��6jyxV�����w�����~bf�R�gu+�xrT̪��ڸ;�q�y�m��'�8����,ށ�8���f�0�ܢ*���Wvݔ��y��r�J2���G�{�2ѵ�t�RG�d@V�C
�������~ .�\�vʜQ=
�9�<#W�ͷ�wΕi��@�lA�M�\��w����w�)
��*��9#ns�wѴ�@����;8����h��<P�h�̏�_)$۱��T����A��y��/y]�r�U�lV�ή��l���� ����k5�?g�}+Ь~����Ě#����N��u�r���p�*$�1�9��AQ�u�;q�Z��ΤJf�a��H��!H�;!�+�l!,mz�JBH`��5��#�F�[f$�ຩ�[�5G�}cG�q��}ȍO���GK��N�䞍p�6ͦtg��<=�{V�K�4m]f! �?@�O��Z�]*$�K�:����А�R0�O()�f��J��_��&�Z�n��Ru�NYf �e�S�`E�Z8��R��,��ǚvDБ������s���O�0)}*���ZV|mC�+;%i�	DJ�)�>I�'L��%�@EI�5�n��a?�\-�/.�jn��]����
�SR=xW�mBO�S������a{�)�è�繑b�
�E�{l�N����[��F����@,����?MkW|P�Ʊ\Kz��������u��"�����(���� ���!�dG'�%��d�2	�0������;���ɴ���"�[5杊�Cc�et{@�#�|��U���n���
Y�'�e��X���V���dT�s:�i�=Ge~�b���h�da-�LB@@��$�ۍ���3�l��S1��J�����T[��1��Ƕ���G�95Șu��X��=c����\�.M��Kx(����Ƅ@|�Pn��k��{�"jX#	��Z(z�K;E� �/�W׵�g�4� ˻U� �L\G/�"*�e�7���QŃ��3}t��jn���˯ħj$�|�ulFG�)��w�E�~������Ex���.��3��w���!�.3�C�~dP�ݗ�������݈/T̷�Bsڠ�U��;�v�&�w��,�Ow�����Ɲ��)����^��p�5�8��*�����Ve=����Q��[徉}1N�7"����`���v�Cs�9z%O�z��F��o��z�R��C�c��a4`{`8nM")���(�l4]��)�'tё)�����\i��Բw��sU�G��,�͊4�Ψ^*l���Ӥ[j�3fG��Ԉ`Ж#�u~YUO�e�P2�d�}摠t|9b�}eʼ���[���7x"D��l�"��wzo~�I'��*�������j�'Hjz������Ӯ�׏"��������<�Ǌ��8�y��u�r�B�}� �<��|��[6{�,J�J�TE?;a�t��� M�v��xɚ�O�3��%����/3���J|f�����շ��(�?&�*�,.-S�w=v���Z���9�,��WG(�^	��A�:ԡ��
�'~ح���fɨp_i
��S��A���H�B�]�쀅�P�jh�d�/���<�`/�
K��v�d���[8e�ζ�J�2�V�/2�0*ɲ����?�I�Q�2S4;;郡��QԻw.8�~�Q�#ץL/��`��%�����h�K���?�'s�'BJX��\�,v��^���۲*��q%k��X�0��>;�ǝ�':������1 �7��8�5ӕ�4�/$!U�&�p�k����JD��5ǚ��&�\Q�?+�^
 QNp֗}EA��R�L�R:<�e�����K�O��2_�t��b�kSl��&�YyF�k�6�P�"Ci�#6fK��r�nb0�F8�o�y{��{_C�pV�$�nRrOd3B�-�
;i��)
$Ԕ�zu(�������3�m��À�c���}B�o�����tLǼ#C4�a��,g�]?yN[]BI�%���?�C��k������"q�Ds�Z?�↶�sU��?�I0h&!܆э�l0r����(VlشQ�AG3nlp�X��H�%0FY�{�̗D���D�I��6ڽ%�F�$��:d��,5M�%�uڵ�uxoBü�l�N������`^��8��5��Hk�]���)D��X��
�ʸ�/��gbL����E�$8����Ô��2�#�_�Mnq�O:�z�Z����!���_�Ro)-I�Z�6������"Bh9hqe�Ѐ`;(g&��%�+�LA�d��
��NfQ/�>�n=��Wyo���Q�Hd��d/>Y�YT�����&�\U�M{)��N�TG�x�$��CK��_�	��$�7T�,�tŹ��=2|�$�!\���Q��3�a��2�l�ݑxq��1�O�_��i3'�ҞR��� ��vZ�����j����'6y���$7�?9�6��NϏ��vD�_�J��L��8)��Y�Ն]h��͍����9tG ]�g�g?�&H>�<@f�rÃ�C��l���Sl�	��r٪��R�^��V�6q|��p���(���<�~/��<E���w�N�c�?����&�2=~��1�HH~���,�������c��K-�W����k�r?k��-CQ��7���O�-y3����e�ְUz�e�ͭ�����^k�]g��h��T�ˡ���ݤ�U*͈l�]��ʌ|�ջ"������+�ϼv�
�(5ϸ��bf�zy�g����l��f�9`|99���w,<�p˅鮃��yO�-��?����
�[$���<��G�-��F��5��ƹ܁���V�%�9�u��f����<Na:�xl��)��H�3� �����nV��T�t4CFT�,�_��+�aE؝%O%�fm���B�ߐ#�0�S}�ҵNXj���J����'�!�q/j�28:l�L�o��sqhP �/I�N�p�r;�:H9B���.�s��^�vz'Q�Ց/	<��S�qp9]"��uĉ	\�[��t���M��8��.w'h�{���6�����-Ո�[�}�Jl�c�8����G��̲�m�A��%Yԡ��.�(v��97z��W��rԖ8,���Ex|���ΥD3��BRB���g	m�	��a<u�c.A5e�Tc�d��H�_ ��8ﺁ�(xj�%#E�(#(�����??�@k�zc��o91L��VnP6���x����`Ӌ=t�	���;iI���������,e$]E�r令��؜�f�J].l+.�c��Ou����Z����+
�\e�V+J	,M���ɣ��bد+��hg �!r�4�@@$Z��Д����`:$���0��ߝ(�Lv���D���(IW:>���R����6�V��|8�wƟ�y�?���  E&�f���>���@�74��}�5(�)شcWx��oAOݝ�}Mh[U��5Go�T&V�eP3���{r�Q�Z4��IѮ���2/���3��B�s�ѷv�,(45�T)*�ݼ*���%k��N8L�@�:�g� /)0�� �0F$�_��+������B�\�뇔Of�4s��J��CB}]�9�#Z��x��uMSv>
S�٨�d�ɽ�~ep����	�i%��Ss���(s^7)��Fz�A��J�&O��;)�\%��j1�N��c��A�6^G����+V/���w6�f�����ؖ�S7�h��-���x�DXѮ_�̀h��K�X��o,)b�@��[��U�A�����qU 	�Ά�{A:##���W"qG�qW�Zf�0��탫���t�;�2�v�3�1빡Tw+[,|���*s���׀n�۬b4�������q��Z� U���k��ᶶީA�&O;2�{�W�`�*�5�Ot��$GU�8u�%�������(%�,=��{3�!U���A���Ǌ2D�(+�^�A�Wq,LBJx=�˹	��/��Rh�  ��Az�"qt$���y�'�C+�}	�E�����~)��:�@����
W�3B���l6����䲫�e4���|�8�h:D��x�ɖA�i�Y��qN�G?Bm!�Y��Z�9��#��>CEMk)��35�ܶu���<'�*Uz;u\E�xd%��AL�
��M�t��o���(��{�- 1'�p��U�˅��s@p��≾� |7a�"�6�����K8pZX2��w���SULD��n����|X�P _'*���Zp�]�C���0y/*����U�K�RAb�7Aw�H��;�oqࣞ�TE;%ةjw����ơz�ePl�������	��jF
m1��ӷts=>������C�� co��2y�6u�{�Y�f�4ZO3A\�rp��M[���-�4�W�/HQB#mS����
�O��!�L�I��0~�=��`#���ɉE����k�[�d�Uˣ�۶y����l}�O�.�|G!!��H*z>�;�V?<��'#�3%�,����F��������)��O��������P��T��A�ZW�D�g�0���p3�h\�"��~�2�e^�$(�Z��@��谌�G��^`>��,7���i���X4琁�p�������Z�w�bYIP8��S�d~:�RЦײ�C.�Ř5��a�'.�Ꭹ�Z���I�+�'��N��-�{��??���J�XK�ݜY	��Fދ�@7� �̎�ݝ-V��������!Q@�cx����%ՔKI�`5?����ml��#(͂�>J���$�34b��\u����%�:�ª������z�����k^�6O#�qr��)�ƘU1G����z�>�Ȑ�k���#�T���8 `����t����9���B"$+��?��n����V��6���M�� >�����p������k��]��	���@d�2]���徹8폝�k���I���{��H���)١��{v#<.���%o�!"4�<��g��g�i�Ob�_K;�!X�d�&%��a�(.�m��g~�33���v�f~�Ie�~ϒ��z>�]��+���z|Y���v.�Ll-9(�P�[�i!a��L�ܬ�*;q���+�8	R^ � '�6�tj���ɾ��,@6H�z`U����I�眫Q�i�e*�c,�A.C�i�>����ӻlt��>�!.�~���;���ȓ��}m�su�SA����+���՘;��tO3���78h��zN;ڀ��v�G�N#���Q�����_˞y���
�V�R��J)�VV���n� fAi�E�re#�!�T�SO���GTu��{��� �_�F�o��KF�����oCj2���l��C�r��#z��������ǜ���*���w6~�6����Ii(�������T&Ȥ@ ��߀.���1C?��e*��M2�2'[�"�y$^�	G�GXɮ��gjB����s�֚��w^�Vj�bZ����Kz�ˢ>)��_Y�Vڠ��7��,��bݜ���<34��3��X��r�x#z
&�YO�^�`L���m��PEtT���AVAz���2]����y�^?�n�Šh�HZ��ݲ�d^`���e�� �U;�L�G�����A �A�Zk"�;�����<�s��� l!��9iry���ke���"�:%�s\Pg[��=2G�^��ϥ�O�<�����kȅo`	��H��)���7��t��(�a�%T����œGFep������y��}}�o����P�0ϓ� s��q�wxVYl��y�$M�D�Rw�ʶ�9�������`p�9᥵)��zM�ЩY*�jq�W�@%*N�1Z���wDC�IFe*��?�n-�,
f���a�Ñz돮�i�y��}��u�ҿִyU
��;�50+1����aA�j���8ٰ����ס`��(^�kv�6��v�?s���������z�w���ߝZqL�M��0�!׮9���>H�y��3������<}�Z����k�0�������SLY�n~�	8��*8Y<r6���B�����i���O���Y��{����M+`T"�N����.�	4��+p�%�q�XbVxO�c#z�6�S�'�l����.�Ӳ6����W��y�I��|I�j�@�;�R^y���s/�?"�@7�c4�I�*{�jze�U���K�����RB��?�ci���e�\�JX����<2��3�3�z�/��u�_�����P^K�ܻ��S�t[�lOK��0>�0y.9{��}����f��?�;~.���Q��'�n�yٴ_��Q�z��l�+@��spī��C��	�Py���'���Ը���?�1o�ٻ�WT=4���M�z�qb�3oհH�UB}�w!�$�9�.��$���jh�8�!z\z��-��Y�;�noR�W`O5G��i�)��to.CHY(��.tb9���3Фx �� u���C�N�Hm���: ;vZr���ښ�}�.����o.6T�w}��������/\�)�U�$$C����rR��HSG)u��~���v�=��$c'H_R��rբ��4�y�����́�O�K�k����Q][<��֯��*����'$Z�c������z�PJ��ц�����;������u��0o/�;� �CY�Gr� �][=������'����ϦԢ���gN��'>��W!j�'�����������(j�n�>�0�rp�D	XSI"c�Su��昋)Fzl7&ͬz��\>�����oa!���O���.ڬ�Ɖ�=v�~�N���Qۊ�|�~����S�=/>��5�11�����to�&=�o��]��09x$��aÝ����*"(�I	A+u�[����\�u�O�����Rm\���'�z ����2W�D�c8}�������6m12���TЉ�!ڹ��6���	0��a�h}�c��DQ9�>ؘYk����|f��k�cbU��l#3�� ����U-��c|<�z\�V,ՏQ� _<P�5��p�. ��!n��ή�S�M��Z��ʤ�P��s�g����ruM�.�Y 8c}�szq�H J%��s�bDھ�1�Zݬw+�=�.���ʅ䴲[��3g��]lf☌�U�A����Ū''&՞��A��&�A��J �F�u�1_jqjFw�����_�A �F!m��>�f5�nP�M�Q�9�:�I���֋��Ǚ��^���$:Qc��sx�i�/t�K��$�A�%N:h&ڴl�ݑ�K�sq���G^��i�A&�4��F�-�8!�uԴ�]uP��?��}��ñ��uu:����$��� r�^@�Q�ScC'��(�>�DS�-�f2�� ��#5<�秺٢0�\��\�U�3b���*U�ٳ8�k&&�Z�"4�Ƈ��.�T]<�]�'�����v��l��l�����71Q��d1B�1�jy؋���+C�!?�׀G򫿪��`�߈-a;� ��}�a%*�g��%0LZ����n�%Y�:��P��,���f�>��o�1�D���jnJ�� �, ���E3ϟf�� ����El�=?�FDڶ��Y_A�A[~��ho?o�Y�b��䋡0���KB��N���[�ޤ���|:w��U{˚2v�O�=�=#$C�l�L 5������C^	���bD K�Ƃ��d����n��G�nW.}���V �Y8�T�����:�|}.��B�[	��߹B$�3�����L�z�K�!���Q1�xǦ�K����J�Q�J�[uv��*�E��-��P���|��	���Y~�o���U#j�9�Go��^5]�w����s�gV��܂-m�o�q"��p[�D�KӾ�����U�r��)��(�K�ɦ�>A�����f�qn�XR.�L9���֐��ڦ�fK��"V�E�to�`i;�¶x�*[l ��C+��G��z�uk8q��[FF;@��^��� `O����th�G�5��W���F�9�;���Ic�S�㽹\�)�x��KҞ��&�T��"�M��8:��f���>���D�U��^��t�ҷ$q{�W|P�f�hE	W���M��h�1n���?��Z����g���ny����l�/���ɍ�k�.u��{\m�3�]�7g�}0%n�;�|��E�a���R�x���L���GJS-lwֺPY�M���G��TkD�/��E�.7��u��M[v	��n)qck��;��-�N�VI
S��i��(���5�n��P5L'�ٻ�H.V8��+�ҿ���;ٌ~dg	+�q�������GΖ'��\>� ,��4]�[f���F��Q/��V�j|@XH��Y�����m����:���9�$C-���O��{4P�kXKr2A�+8��=s�i&QX�׶a0�h	6TF��@s�;.��r�k������ѣZ�Y.��*�E���}i��!O�(I5�Ng��	���?��&����6�F�]۳��	Z	Ud�mu�N��5�m�EO��l��r���-��E�l��Ě��i�9������K�gW�V�մCFw~=J�*"�]wf��っ�YV�q�֌"�ߖ&(��4��O�;-�B)݌9��{�ܞZ�6=m	�%��49^�6�5��P��9+�5p����B����mϵ��P��9�/c/�2������A�9\����n�� ��'v�j�&d|�@�X��2М�[�=�C�����{'��Хh`Ķ�U�x����Z�E��7�c��tyaz�L<MnS�vD�"��#�.�jko��N�嫑�'�����h����/z���/��"���Tx5�wI�d�QHhtl���b�Q��|�E�Y�}ò�?�C���\���C~��;�/�4c�	OPA�9J]��*�a��j���.��L�j$�0�uзC��*���>i� \�bdwȨ�qu'9q���Y��;���>��"�u�I�w�^%O�7?On0��e�G�����O�@�
 �]�wyn���K���O~�.���أ�l�'JB��am�`P����kǨ��D �K� ��?�I�&�����"�+ݷ��OPm��Ū����!��BR4����aa,;N��{�dPΘ��o4['$������[:����HG���_o%*����[�CK]:�5|p�q�����l��1�"�=�M\��A��o'�Z<u]�1�?x7˚F;���dP�� �a$g�v�3���JI�ӭ�c��"�u��Ytʫ�p,��(���޽F^���c~H#����z�@}ҭ�KtCh*�O3Ļ��$Q�7f��>��v�9L|�말��*�O�`]
�ohn���X7��+<����rGΈ��ﲒ����3����㮶5r�A��ofk�IQk!��]x�T�|�ͼ�(��u{�P��#���*�LT���J	pŧ���Uy�P����=΅�=�P�6�����dv ��v5�AWj��l$�u�a\a���"�C��jW�(�W��ߏ{<Jܝ̺)���U��'81X*!9�9��V��췃h�c{[���8M�����K��(��,��7����F^�����{���LOh`g�N
d��� ���5��|�%��c�1�G���?c�'+�Pi!h1KG4��y���w ���P����E�Q�����N�J"�C:�[���& izZ���gj�9�"ڳ�@�g'f��D�`�^e�/��(�ȝ���}b5&��q��RL	8�u�.�o�{��">L����	�n¨�,���C�"Қ��s{H�3kc�s�j�Z-[	P�������2~�l�L8jߐ��u��+F�� �O?����w�� S�\~����d�C>��������|P��
F��԰|Q
��h{�o�13^�@iPY�� �s�W�y�S���wȜ?2�{��Q]�P�Pؠ��@�BU,\P�xu֓�eD>���[^�,�Lv�oJ >H{CS��xR�z���v��ݿ�r�j�- OvBcX��	�0?��W�z�����m@srɪ�I�M��G��o�]��k�eQy2�����:5^��t��j�6b��m7�F��3�%�1)����E��}/�/r"�/H���9�.�Ϸ�`9�ǖGɆl�����h���%���z�KR�Pa�(D��|�N�XK��? +(`�2E��ei��{��5N(�%p��q9Nx���\�J$义��^b������3�E|���xU����h��{t� ZD�K���e�S�i�Ny��u:�/�����3�{-�q��R^�Ӷ��FY3�q6f�/2t�3+\���%�`�<�J�"��ҩ�?����P3dt����ŏM�h�����X=��S���Pp��u=��$���7������T�]ҫ��!m�ЫC&1t���F:Mr_K��(�],��v����D!��ܻ�Z�Z͇��$���Ѭ;%ԯ�j�E�8`$���u�}^IW�����cZ{�����˕�Vk���^�	煮+��LI1[�fRR2Y!�ޓZa*�"[�F��'���k�+�Fמ�44��D`�Z3�l5? eÐ.F��t�A-��l�eN��{�d)�`� <\,5�������Eg�XO��.	���[���Zc�1Ù�eX@`�[��K|Vam���Dk�ӪZ���Հ��AkL�p�^�"���������f.��Ew�m`gr��tF9�ݚ���e�J����$W�'��j.�����.Ω�/��Ĝ�����W3+�4�U�W��·�F�FWG�"����EL���_o
��b%2�q$*Ux�;ޛ�\P+R��~.Ҋ4lV�Ո�v\��'�a���b-�6<Փ>�����u���)D��<���]��/���K�Iۥ��O�h��whT����ԑ����������45��Z�!�]���##�82=[��Z������x���%��W��GAy�u�p�3�����]�Ľڄ���#`�c��^e3�.r�ۼ#�<�o�r�h�Y�(b���l�v*��Zi����u�-iP0�sw\��0�E�j�8����9��oH�쭢�N%��mAT���Cm�� #�����R0����x�Sg	4�G�/4��)��Bg|	�g��T��B�sI_���`���q���Kk��1\��{REnC����a�B�V+�IAZ�N?��'L �dG���RX@M@�#I(?r�Dp�EI�G�*?Nh�oq^�L����N�'F ���tv��J&13"Ŧ�OD����PD�Oa�R�}�B���js3��=���p��h^E�gr��'O��?V�{3��ޏ��Z�/y��i���p�H�B�J��H_�W#�t)q�
]p)&C�?y�=�{�R�LFH.8��1p�6�/:�X�6���%� �-La�1�N��t�
�@���k������h�l$�2|�� d� P�
3�F-��?���C��[���p�3�L�"��H�FiiX\���eX���\���Z�{����^��fL=C�=&U0ܲ4��(��9JVB�-D�#i��'I�Ю�>������f�!N��E�.gk��,�&}�Ah�O�5�JbT �T_�C5K/g$ d��������
�@���%����;���7B�4��+`%`f+��d�ʀ%�&=���$�\����>ak �h�Ȏ�^�)���1!��� ?R�Ǫ��P¢!͘�*��M8s���gw���z�z��X��مP\\��}�]����!�:�[t��f��('���B�6�!m�r�څ��N#��S�f�d��i@��w�����h[h]o���+�c�&lG�b�p"A,v�����V�������&cֺ�1)�����Y�p���Vz�lڣ��U,J8�����P�1��-|�4�a�\�����5�m�,��=�}�v���P59�oK2h[�#�T��^�-�UǍ\3����v�y�K�(��%�_�D����H����3�������ȷ�����W����n��D�����d���q�Ԃq��qu&9
�����&(�`���
�ZO�K<�\�
��.`"�搽��x���`-�+y{��h���y��P�͍����;�O�w����ݿ��D�I��c[�X��'�{��A���/Wp!��{U�H�HH�<(	Ϛ�`V�M�Aݚ�[e�ig~|��"#{�]gT�M�K�\�%�m����!\K�Z����m�б��M�s ��K@R*�N��e^;i"�D�4߉�C�9󼼽�����5I��`�U��ŹΈ,ћ�y�$�K(G�����4�Ih�NP�e���QW�����-����w^���/U!����q�G?T5�m���v���I���;��;|�*�Ub+��
�n�r|�=q�>EG�hi�J}�b}���V��2K������A�mT�bx)�n�'�ڹzʛև:�$|*:�p)#�i�(s���#���e?S�b�T��RI]��(?fAX�ߧ~XÝ����y�Eze�g�)���L���j�LB p�Q'/*�L�x3� �DK������*�}Z���Ğ�#N�JT���Y��ȵ��K�����:���Ƥa"�/�L'ud������i�b�V` XC�����opD��
��t���jh	��:���՚vk�ܿt7�-�e�ȡ����wb|�O���|B/��<|.������ɏ0���.i�_H*&\NU9�~��=t��� ��S��$�ۄ���9�����7��Ҡ��4vRa9���۝��0.���W�-��r��O�*��a�����D���O���@��nqg�pQV�s�^p�� '�
�����.i���/�E�ˣ��|��̗NJ�S�q���fs�!J�����0���"�c����������l$!�aEv/V+\��ڮ�V�G?!n�/��ZV�t$CD:e��7�U�ל��pi�u8�mp��lZ���E��4Ķ�C%Ӏ�E0�����C�j��a���(�>��<�&q�O(�=�B�k�$a<����P�MMp�) x��<�.�>>�[�Q�����i+�R"�S�>�)^���ƫ�Y8�ۏGBu�VI�U��U���?��h�Q2'f�^ՠ�0i����._À�"���(*pL6�B�ߚ��"ZQ��仟?�8��FZ�Fϛ�&I`��6�+����Xb�p#��Z7��N�_d��5�Ͳoʿ�4�I2��2	��ǟ����3Շ�Rb�ׄ}B���|$3l�^����P�,�IO����>�m��}��K�ၠv�/�zi3P�j�\��p�X���u�JCOZ�הL�fw��%*6����z6���y�S�q�\�pKd�bd8��ҵ%I�}sja��K�xǭ��w�2�`}+��w�>꼑����wiG�O9���g(|\�<h+!��g�ٶ�;MS����h��<�ya�����%�;��r��-�LX;uʵm)3�6��p(�p#��U֦�d+�H��O{�v\��É��;e"��_����渾�����H>=!K�kC�}K�#�j��G�o�y�Fj�W�#��#��2�����l;�/J��i>��׻L<������Y*��s�@����%�ߤ:R�8��[��M0�	1]�C��R��ש��wV5N[��6�V��cv"�Zw�B�-�w&�2$WU#��hVϢ\* g�]���iZxE��.����]�����N�&� � {�����X��A���ٝ�T���󫎘M�fn�)h�W��fѭo�G|h���Eu�39Q?�jQ���Uh��3$���᧽�!��[�^4Hr�iH��T���Uc�;�h�'K����'C�c�	&�t��BV�!=&��I�v��ӥ�����S9�.�I�%Z}9�}.]i둾d��Z3��f�r[Cs=$k�<➥�3T����҄�M�h&=F�>߫B_h/׸uM;��>��@�:��Q�0���@��,o��)��SJ��t�<f�a����u�1�*�@�q�'Շf����"�B�@�쪫y �m 2�������ss���C�oţL	+�Z���V��������^zd@vw5�s^Q|֛�~���S���YITʹ�?S�E�m��b�7�D��>w-W�ҪU4���_�0���1� 0Z3�c���}��a��:�my�	�-9U?R(;C�d���eK;����y�+���c�L%.����l�`K�o/�0�2-�r�M���Z�B=m�m�hQ��+���tŜ�ו���r���HHd'} ���2�Y� (+��4�19�؛��%g��lʽ]�,Q-���^�r�I`!��������/<��!ԫ���h�{g��\�F!�͂���=Ɖeo�dg���!�		',�~E҈EP]����hX�����D6mo~��ܔ	 �n��9?��.�GW.K�S{��ʎ�X��z��`�3ٷ����Kfa��Q�nQ��jt�K
��H|5�'T�#��bOx���7Quc�.���#?DvL@����֢e��A��(��ш-r8���Zՙ�ȁsv��3.m]�z�=v�N�mf��۲_���t+~�(Y�l�e���-��IU0��_����WNJ.9���o���F�GI�Cډ�d}@~����NK$�n�տ���i3�jo9�	�B�;�2l�Z���q���F��#V����6���k���rr�z��g_��Q3&����X�C"+��&w͘l#0�͕�r�h����w�uh9��sTڜ�'�����*,�F𒧢��R����m��3�2�P�RBz� �z8�HT~�1
�X_�	��6HI�{���g׉��t|��:���-����T�S�2��j�I�ORː�K1�Ɓ���6% 1>.��a[�mX���0W��T���K��1�鞾T��r]yx�*�ם� G�o���od�j	p���Z4kc���~�FV��u�u�KB��2�� ��Ek8��_��R��[$<+9�ʅ�}��ՙ�^Xͤ���}H���D�����e���[1���OT-��������k��J����A9�5�������+���*���|#�!��ḋX�����2c�J)��Rrq���Yρ}�B���W�����EuV̔���C�����R���&;�\5�0�W�V�����r�C��
s�SP���ܝXNCS�iW\ܺo0x�
tO��
����JN���� ƽ��6�d��dE )�:���}��p��D;[_�G��oUE������R��z�
8�?�	%�XW���uE42K����IYחx�x� ��(�^QAq���k����n�J����� 
[�� �q��B�
pk�m���o�Yf@^Z�v}�<v8�<9����DQ�R!�F5��'�C�u��G]�q6�gE�׍q��w/r�ػ��yG��B=?&$A���91%�J�^K��z͝	���Y7����z����X�G�@5۴H�/�+�ۮQ
�O�^�>�����X��9���8�*�Ǧ�iy�O��M]��wq�nRc���U�{��$��x#���yA���{'8CyZ�{0�A;ѐv�;{����_h��K͈�ނ�^���z	��H$��L��DD�m,	�Y�P���X'B9򗵵=� �G�ӄ�܎�K#�$D��=���/�t�2�|�{ix1��>�u��w h?�����!�+M��&|����ڴDBJ}����������l�&ZW���4W,�RK+���P���z^�!uE=��J��S{/�
K��"ݲY�F��/��?��㡱�R����+:3��2�s��ֈ��� \�0l�ͩ��֓�C�������Ŭ�>3��Ji���{(ea���t�{4��Kаt�P�|[5�%�% �	����Wd�5�*
��6�K�;��sM� ��FN<�C��v��T���@877ϮI��iK��ݭ�f/E!z��qo�T/�7��D`���a4{Q1ڢB��k��R:G�0嵪%H`��i3�B�E!�?d��4�A(u���'��hzηܠd;EPf��|��&�v�n�o�̊�M�k�f���"�3�n?0M��ҍ���@�cX)n/��(�\C��Uq7�1%'F�og���d�7~��%��q�<WO��0��\YR�-|��k�p���jDy˄��1n���ĵNH�`�FYo��b����"�ޘ$
�@���M�.�%�в����ʴ����x�����&Х�d)���c��0r���	ٰ|�A���*[qXR��ߙ�B�5z���䓰�j}�v"�
Ul�ð�4ꋇp��%R�0���+�$��*��&��KI�c�,�3�5r�2E*����F4�C�=[V�� ǚ�`�^��.@Z�<�x��^Dv�H�Q,��iY6z��ׁ��#Ɲ��(p��חa��ŴR��"��V2���¡{P�e0�b�;#F�e�x$d�}R5"5�b�b�m��b8F���
}����:~�4æ�w��G���=>��������;��ƈ3�sr�kp��J���}��,�3;����Ơ�6�M��-���\g�1A:��]X$�F9��ꛋq�T�Y�J��H�����>S�0��֥.�\1���/�z13uLyƘ�B~�T��o�5�p5��<Y�FC��t�]SEQ��W���Dn \-���/r�8��J�H�Qp]&)���]_@:��6q�A|L܆B�4J8�K��R�m���ꇤ����(�y� �t^��7�����V�����@n�Ǚ��9�yTzG#�H�����E9n�Ja��\2������&*��T�T�\��9��t��-�f��;� �J��sȵ�rv��6Od<�R�Y� 7� ��UuΏ~��ڴ���[�����g���ZBp�[y�I5[�����<��r$�!�i����B��A%L(�|�H���I�Q�����g~�#}7ǿ	���W�ҡ
�"R�Yo�7�)���y�|�8I;���A���õOB7~��~&��m�i��͂��QupvK9W%�p�q%#�/�f����`
pPH�Kg�����<m��4��I�ry��M���m̬ם�)-l���b�	d�a�:�45uB�x10k�U�T�hvH���T=b��(�!�`�޺�#�\&E�ф��r����"M�`=5���_��5r�?��u;9�Ep�y���*��Q�(�I���B �)5����j5���G�������h�:�.��HI)M�� p��pO$^�П���T�R��\�<�;����<��]�n���[�hjN�a�D��eg�c���XS