��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�\a��YV4�|�2�xrg�����<5����ߵOf=���GfE�����ŔM:2���PF,����7��7�� 8dX���e��)�Ÿ�k�[�t���Ӽg9�(�i,j+`�W���Gv�U"λ�(A|f�ﮥ�&��T���T�q�CJzXu?��3Okl�̋/��.f���W�Ė�p��')?�	4��j� *ܸ!m�q]�Z�wuعG6���,�Zcf$�]=�����H�������0����=��9� �Xp�?��)v�� �E�ﯘd�����`E�֢�.�x�:��K<���|gL�z��	y�d-���|�ZP�B1��������M�Qv�Qz�Wơ8����S�� �60���P��5��$2`�<�R�  
���4�U�CA0�/i�6�d�}�'�s� �L�.��N���|$�qyՙ�B�m�2��(��ny-�P��k�%�g�X/�e��Ky!P�P��(L��-n)��{�{��T �Y{�|CK�Z�?�'&2���Bi�i\@��]ix���l��d�X�럽��7�IE�O�BRJ�K�������?���C��M���OV����Ӱ��>�Z5����J&q�o����|7�G4Z��񯽗��A[���8+r�b�Z�\w�#��E C��+s��6�n����B?h�?+ް{�iv�(J�:\��察B��S��rmb������=,��U4��`�&'�[�z8~�g5��9�Q��\g�d5�/�뒕V���<Mn�7	@�ĿF15x"^�r(YtM�_�Ԁ��D"��%^�O9��8 en�p�"���iM�'R�H�+�e|!�MV,J�4) �	�L��
m�Z|��w�Ϯj����36��EB����q�%����6A=�/��K��5���o>{aE�wk��f��w{�م���Ț"M��d��0GA��M��_���Z��>K���bKƬ�}fq����(':Wn,�8�J��d��ڸ֊���3v�t�$�壙bl�l��,�U�w��<X,�+�V���Ė-;v�D��or����Ɛo)F�J����P��1��C��o�1.9�^� �]��S�;Yj%^u������
��A���j��Q�a�6��1e�:�]�O�ؗ�6��P�3�K|j�sW��1����y_���4�q��U� -�����-�K�"��PW*9�~q�XO�M�������f���~��=���@�p���TR��=�_Lÿ��jv���)�߯cA6q��Y��^�ډy�h��i�~�V�؂�nm�M�Q��7?1�ݮe�r������M���`���T&��F�ZFwp�~۩��lC[�]˪��)� ���#|F��軛/|Wsk6�C��ž#����#z�H4�J�i���nfV��Kbϸ۠���y�*p���W@}G!�R�Kx_�W�'O��Ṻ��;s���3O��/Ҙ�� ��\�}�/@��zR���P��	�(�� |��'�:0� ��9�k'*����z�h�� Y3�;��ah������N�/mʞ���4�Fq`�s~�b�/�\��oJ\�j���$]�g��K���o�"G��.=!v�e��h��!���6���hu��¸�ưM8�j�@�Bͫ���L�=���ы���3�9�	>�k;-+1�\�0AB1�$\��檀�����.*\͢Lؾ-��r�-��`�;��=V����o�C�� �;��Cg��Ŕ��I\3����q�>��*��Ԑ��shlh��*cI��B������7�ՙx�m��E��j��g��,��	�%u�y iBz�Rݸ��xl]��[�!��`����3�~�����)�A�j�\Jڰ�s)Rˍ�Í�� ��d�d1�����j���� ���+ʕ��Ɩ����>ʾ�6*���w���e^������8�Z>�n���qwm9�5f�_$�X�G.�T	mFs��}T (���|uaj��6��7C<@���I�:�(�o~L?C�.1��-d�ś�Si�n��F�Jzj�b��N �6�Y�H�E�U��B(����C�l�8���|�?���Н΃�~IA&���Id�,��}��y3�#�R�VѬ'V��w�\f��FN�ƚ q�9"�1���Q��Z�6|�����Eѕb?����I�_zB,��ݵ�G�Ik62��s+�izp�8�P�^wU0W���e���~^Ia����[qK���u%�f��U1� &zM/۠wA±!3��I(���J��yӡO���3(v�s�v�}�]*�ʔF�ڹ�'���\W{���R��`V�=lLP�oC�A���("90��ɕ%�X5�:X��,��}�t������Q�S�dz`��|��/S-�L�7��`>!`�#����J{�N��"fh���gKG�aX�"u���V��Sbp�n���J+u<��~�'�7aS�Vb�����(�(W��j� �҆g+�&�Jg�%�%0+j�x ��J��m��M�Ě� h���{o��,��{fܜ~Fa6
��Q��;�Fȟ��#�����(�ыH��;�U��1�l�Ԝu7R�k����͂�_����=Y�)ɤP̋*�/����I��d���
�K������ў�L�Xr1K�N�R>���I#�z�z_�ceB��^���*�:�D�qsFa����&��̿+S��[�(��4�{6��q����e��R�Ë�nG��!w+��~�/;CY��6��2��|��j&���C�Bu�u,�d'���P��+�T�ۖ����U�?��B;�P�tѨ���u�;��ՐGЇu&fK'l�����Y�J�#��Z��Wӹ���(. �*�4����d-g�*�t��wI�;�����f��.���ſ��0w�L2<ܣCk�&��e��g��R�r��l�Q��
�Yl��3gW�h��������D W$^e;��67P����g�_�ijfH��#��MȊ�ɷ��A��&�qH�5XU��2 [��Kv�f�L7@�*j'w�3��ކ�+�2]�̦U�n�e�?��O��w
9>͠d�酴�s�FpC���Ɠ�c�C��f� �R�nV�W�נ
��xdb~���v�d_�(��Ț�X�3J�S���ֺ0O���mnX/,��Ps���j�%m�}c����Z���7T�5&`P�@?��iy��YM�ߠ��}[a�`��@Q�P2��'慆Ep'l�n�75��E����^r{[������AAw����<�1Gnu!W�ޱ����e%pq�89�f{+����g�cT����q���ǜ��.�^>�j�\�w�
'עe��ж%eU�������o�][��� �/��j�I�s��G�s%q�zU��́�I):�R7ƕ����/��ǂfA#6FH�_��?f�G�Z,m�ռw�{�gߒ�����������a.u��qġj%@}	v�t��+�t���{�����V�X�,���Qi�i�}Z�L�t]\��]Id���p��
��2�}��O�����J$��[b�lu�������K~�x5���%*�I�#u�y$ds��p��=B��:�}`{��<�,�H�o,���F1��k��O6*`�=it�6�F2GJ��s��':����Ue,�y�=�xc^73�Qp!�r����N+.T��]1����q�m*� �\:��I��̲���v�+�(6W�[Թ,�h�V9�����%&#cx�WB�z��� ���|�/���:چQGWV��*U	I�m)g�E���u��Y[�[艤7ޖԃ�E����&g�Ϡ�� H�5���dH�h�n���^р�˂sk���޲�VY�d�2څ_�Tj�y�n�PL<����Kv3W�ߡ�y�.��dgy�r���U�r��T�*j$���kV������iJ݁���ܑ�^	tJ�w��l-��WWp��1�/�I57�'� =�Q0-�[��2-a}-<PT?Z��q�.g��Fx�vz��M=�)�*>aA	��)���[+�� ��=����:Å�&��t�U7>�Q�]��c/: �D6�r�;Q �L��bD�S��Nό1�J>�,,��P i���?�4pk����'��~�����86j��������@L����%��T��&��nR�ۓ4�;s:�|%�P��tǯѺ̂䍇�V�rm0�t�z�k��O��(<��c�3�Cl�<C!XV49Q�<z��5�q^���Ɓ�&��[����B\�-�/;�G	�E�V-P�dY��^)/=yR����X�5��l�KdS��k�b��e�2�ȹi�m� �t��b�K1����qe��mn�f��Ci�u�y�L?k�]� �  �mS��n�GbvE�f,����D��@�_�Z�2�a(Y�]�8\Ye� g�e��#p��{�9/႖8���R�"��RI/S���mE�D�aYC��L?�ִ���+\���<;a�I����!Z w9�{
��4w<��`�<v� ͈Z����P�b9n�L�!��ׂ<.9�������2���5h�����S��ӷC| ���>���-�껜Y9V��0"�f28���m��Y�"n)���^�+t� 1F�=d�xS����}�R�xAF�"oi�cV���f��s��mȝ�5��[4~.T�X�6D���If�i
0���ևp��ؿ̀g�ŋ�\ME�,��1� te�%��e%q�A�b�g�Z���y�����Rm�[�_�\p��S�H%�fR����`��_���B�v7Ax�ͷ?�����$��ʉy*)8AP�E�PbԚ6*&��Fkp�����c���/�(J5�����	Y��v��y+A�s�A>׺=�_��;��W}�ej�{��-��sI�6\��S�G�1�4�1�\�>��g7�{al��kQ	�������*qXp��T]��͋Բ�1���ع)���� ؒ1���Ò�=cT�}���4$al2t4���=�&�c}˿� q���s�jM�A2W%�ma*����cV3l�VF�?Hl��/��E�*!D��EK�`UhDx�Gȸ*�3�;-���5�T��#��ٷͬ[�B޲�\��=����	�}����s�mRZ�oSt�T��4��~A0,�Q�j�g�J���V�^#pR�c�*���0q�mp1����c�^m�2����ڏ�,o�֜q�0�����ؚ��)��}��d8]��vGAh��Аm� 9	�o����>M��S�9�v&�E��Y�Ā��0�g���ݒ��<V�dx��i��Mw�ph����E��PѪe[�l��淺S73����Z��ߧB̪G�a�rCKp �0��71��aK�l�8�.������_�=��m��I�o��z�>3�|�f�	�yB��U����{mSP,�=�9u�����V̭Ȑ�Z���������&t�#W*2^ʼ�{i
L�d?�~��xfR�Ȳ| ��B�[����o� S�	�џ�A�,sD(���@ �C�12=m�0vT膢�A}��{�ɔ����c���5�Xҡ������:�``��Ndx ��z����P�rȴx	d1 U0��F7�*��Bjɜ���<�x��#n�#�Q���Q����h�t��G��,`���NKǎ��`�H�[-��[Y0���������}aK�Z�P�Sk�u�g��ɰ.�=���)G��ljTĻ�|��Mp��#�q��9*l#)Z���X�mڵ�gl��Sq��S�O��w	J��vVưj�����G�Ukc��$i2l��G�b�$�����e�ޑ�/hE7z���<�L~:�9�R�K��vg�'!ٲ�S=�r˨>j��������H`H�p��A}��n�H���<O#�p��+�ُ�7#4�^�f�����P|��덻��ڗ�f�pfg?��&z/e+�J5��|�&q"JTq�W�� �����)�	(S4�y4��l6l�#:2��]y1{�⨰PT���!�ȇ=��������m��/��!@DB�B��3��_*���.�#:VX���[}���!��ԛ������;�4�=�v��!�&�������\�J��4}࢈��%~�vԌ�{����v"��R�I*����ix�a1�;�{�H>�X�ݞ���,�k~��o��|C$�I@����Р��R�y_CȰ�G����v��:��=�e�Rw2���^q׹|�`�2u�`�:�����Bc��Nd����][�����������y���$��{T"���14�
Z��o�}���(Q�����Ҳ�6 �F�Y�/�]�1(�Pg"
�(��q��2T\�w���/�Fĕ�ٞ/e���|�\\�`�#�M�I�ε|��yS�jP����Q�h	���[��E�YMG��#�J:����P��Y�� ��=�2��"�^���,��v�� Ǿԋ��s��!b�]��@���vaɸ��!g�a�mQ�c��[AC��;��}W�~�ql.8 �p�{Y��խ��
MP	��OU��O�K���_���ܻ��P��	8��HPb�	�=m#�#2�?�ӑ���������T8�O�-�ĸl���s��T7t����f.���姅�pїZ�~?ĕ�S:Օ�;x]"C�v����� �IC�[ �������Y�� ���؜�ߢ�5���U͐wo�D7J]r;4�v�nF� _�1�xr����??�N�\5z��Hy��>����!�`g�#a2�`� � �:&���09[GN�_E&�-����@�6���Pho_���?�o��;f�����a[����t`x.,�N�/<NG�Z#B6�?�ν&�qI}{�O�[��ƥ�@sv��o����aM�Z�͙�t��sj6wfr q���s�X�L����]��k����V��H�4dI���"Y����:����J�^`�w/����.\��>{�Ml
T�ۜ����3��%,�'>6˭_��T��fHē��iY����R÷�یQ_r�B�}X�ms���*!��F���V6Z\�X�T��^Q�vɣ[9�x�Q�k>,lw�������O],�*�⿀W)�(@�W���q)���cq-nؑx��V^���a�k[1�C#�̓��P����Y/�3A���ҥ5����r�?P��
�t��#H ��1��1��I6���\lh
�����'t���c�6� Qb���\$�P|I��d"���&�YWiS�h�W��q�t�������QU�Y��oq-�����H�P��`��1j����"e/��ǭ��3T o#Q�C�<]���]�G|���3�P�
�r��`A���6�Uw��C���_��?��J�4��GP�b���2��/�|l��9�_Ӕ��8J6*��y��X��K$�U�{�x�\��_�'Tg����jag=T���fy�=��"k[p�>\^�U㺺j�R8��!�u�������q4oe����̦�BZj�7M���j/�<��DŖ��X��(G��1#̰;���<Q.y�5�]�*RЄY]��� c(/p�2�ʣC.U���-�~�5X}���e��w'�P$!�h\�"�������P�����ӷ����-}cM� 0��X��l%�܎�V�c�i&X����45��o	����I�����Q�}�`��"pV��
�BhX��'��y�-�YP.^���~�ت׷� D�f� �.>T*�;Py�][����=ت�H$��(����hT509g�v�T��vX�r`*��G)�6�oܞz�rb�v,�E�ݨ��"��G�+��������S�):7OwB~�����q�ݚ��I�3Wp����R�=?��>��ӣ��Ao��T�S=�M�D%�
Dp?���~JR�[�Ya-ש*P�R$V�&�C��ȥ�4]&y�b��K�m�x�$B|�Gs���I���,�K)2Pq�C=��������k���-�>�� l_U��g�ż2�z$H�ZN���I�u�&��F0�1FH�}���UNf�4a����9�9�5�		w���s���]�'J����U�fM��Mm4�(l��qPq2�V*���T�<��4I�t�']n�-`���<���%��Y�+�x��=ǭ�58>\�z@=�&cS<���G��%�1TLR>ְ6}Q������������*.3��Q�6�營�iCR�.����rwW�������v��y7P�sY�k"���~��s0�Q=)?�y׍�� �C�C�����0�	�d�Q`� =p\>��o(�*�A���i�Vy}J�C���$ZB_\�Ȓ߂Ɂ�l�Y�����HZ��M�K���?3��y!ǘm����^C��~g��c����.I�e'W�lL��ָ�L��˹a��T���O26����e>��7������û� *u�a��V��:%��̲|��,�˥$�?��<�f"k�#=�# ���`�}�Fl��&y�=�^k��(�j*#%��-�U@V��i�G��b}���Z���s�R����� {��	%�1��m��{�紆ЍD��a+��G��͟G�(�86O��y��O����s1^�Ueq/Lӕ�]U�&�(}�ֻ�6���PH����-���r��!�70�1��?�&�Ǆo'�s����,���D�J�s��cuN[v�1h��A��nF-&�v��|L�Ol˃#�Z�Q#K��2� jO&~��Zk�n�2Si�Y�<M<%�A���qv�C' *#�3�&��;�Oupy��У�^�i��NYB���B	�	*�׸��x�OB�j��h��5{��(�i��S�sp��c5�?��(ϭBh7w��,�"��v�C���M��	9�M���|��8ӗ�S���3.7W��q���[�L��mhwP��6o;%��>{��0ݎ?S��	�����}籫
��mΪ�޹��}(wf���LY�_HS�F��g��t�ͨRq[>��L������e��+j����B��jj������Δ�3+�V��y*�r��u0�?�/6�����+?���<�vF���ᒴ�t3�S?��;�6��L�\p�=>��#[�Q��9��ͽ<��O����"O��T�#���Zy�ʮ�HU�|���Ŵ@n3z�1�e�2���0�mْ��<.�~�_���Ww�!���#8�3D��]4��P�
es�Q=����`u��Z�=.�:D(�w���U4���-�7�_ݸ�H�EO��C�.��薍p��-��-�K�SH�&fQ뵙��>�I�X}[�?&Z/ђ�m�e��Z������oQ���;���Ą珠f]y��/TV��BN͑�����Q{��2tx^���%A5J��n[�%�zL*�o�����+���Ԅ�I �Ϣ�'����ht��	a4�*d3y$��������x�H��
$ި�����)u�y*���+��&GcF#�i�g�����n L���ƚ|a��E����]8�9����p�][���M>���yR��n�<F���
��[v�Y���֐rʗ�s҆+��@��N��[���F.���~����GN���J�Yi;H��j����T�J�����,)���5Ҷ���_�F`6�z�uy��`��]@�v�b�m�$��_����7퇭2�#r�2� �`����ɮ��̊���YDWvF��-��?��/F5���㑙���r�l�>� �ӏY,��8�2��5{MV�������0�:��2U�V��\g���sR.���.(��z�)�3ߟ?�)�,��o_[[i��W
uĵ7��Bh�/S�Ē�981��ZU���G��k�,�o�ES�:�U�}'�|��g�*p��>.3���0d�Wj�%�����
��K���)r��Ǩ�����;K��u�+jX���Ԗ�[lȑ'R��H�����)�IVj�05.���Z�H| ~���ڻ���B�ϰf�9��%���$=t�3e6_W�jF;=��ΰ�O0�b���I��J�+�2W�``���{�g}N$��9��6��0��f��uS��~�i-���ƪy��v2��L]u~� $���]5yq1m��䲠���O���8c�^)ܣ��R���{-���}�a��3��I������Rrzۚ%#�d$���J-�K��k1{Fj&[�ǥ붯W��3i��8t|����O���f���^�x�nf��Ci��0 �*�|d;�����2m�^<�f6CM�C"�b5���������6�R�8�����ڊ�UMжJ��MU��[f��>A9�d_�o��둼B?⛛�uu���&�py��\0���ߌ�`ic .jc	!6�8��g��!Ӈ��Yj�S�>�{���`�6qQTzI��������s@L�L+�"�N����h
�\ y�G��I �h�����Mf^�R��kBݰ��j�{q�8�A�u��m tfp�$W8:��fC_��<0=G��j�Ǔ.�� ׷-)�9�Le+`�``���R������a��,;�4��̤{-3{KQ���m+n�''�Ί����#_Z�}�����oԚ�.�tm&�~���C٣�I$~�}�8�7�.V����4+�D�$���$~`���x��6(���\�`o�="�؏�gS���ÍE�����c]�T��F��vH߆1����R�oH��fOԓ=��$F_h%�%�z�?Y?ItXd�R!C[�����ݬ-(�87n����o���Bόbp�r�ٕ:�Ae����0n�$�C>���`Z�h�fO�
�|q1��G7k�*�6�N�1���q���f��ٛ�!E<
��q~������8�ӭ,��d���盢�||�b1ޤ%��������	�JLq���C/[R���n�hqM����c��#��S��!g�������v �Ҿ��Öd�Ï6�*ሽ�ٲ9�|��ө����d��
C���'P&�H�K�l[{�
eջo۠���E$����/��=�Ra����nh�wɩ$�$�����-P7�j���7|�I�X�|�q˶D�Ͽ?��Z\6#�-8��n�L.?��:>r~k����/��X�M�˱������q1���3H�����p$?39D�#<hH��{��F�ݖ������%��ŋ���8�.��P4���S��[�DUP�R2��:Q�*}�+a��0��%�}��C��e?"���EE12�ҥ<�����{P����\����:1M�d-�vR�b�q�BKx�w�7��2yhz��]lx�b� 2[�i����cP��y6�S�|%�1��@7� �	a��D�#���������V�*p��IȼT�ĉFiO�`#>���M�GH��{Pe�Ќ���]�J���)u��ՍC<��3�˽�d�����"ה)����� 4�$�����4Qx����k@ʻw���?�%0Uc�a"&���sj�H�y_,�����ф�$�+jR��6� ��|
���(��1{�1D���L�u�=�|>:K��0�,ퟲnfU����'�8���p6��&x~�^��ׯ� �ѧ�bග�7+XJ�On�H<k��_&'��y$
/t|¦f���{�u��\mk�F�Fķ�.�ӊ�P�%����(��+f�G�J,a~ȉ�AJ������Ex���Y������W�(��"�̟�F�ۼ��y�t�z�)�e��VrJ-������k�G�\m�T�ǉ����������a�W�΄T[���1/b��/1�l���R��S�򊿮�&���Հ�ù�7i���F8ABj=�
�}p���"�ئ񍬲HE�?ƪ�]��OK��F((i<��3�"�S�&5V���9�=M���$�Q��&)� ��G{�\[9g)GD�N�"sA���'?y~�NQ�Zw5��f�#��e�&(�o�g�t�yL�����r-�%}*�N*U)��,��5o����[�u���of�A�G�5��:�_W��Ig�ot<p��F3_��w�!w跋
�S�p6\boE"��fU�bo�`�M� �[c�K�Uy�X� =!�72�hL��v��O�gD�0C��ʝ-�oFU���$�]�	��9�����҉.�=�4{��˰�&Ϣ[\���2NN�(�!}!���'7�y̕�!!�t������ۿ��{�]8��7b�����0�GI��4��������Fk��"��Ȥ�^u�aZN��+��,Nl<S���y	}������3�*�[_V��Bk�K�s��_F��]�ε�vI�������l�EB����~�P�4��z��(���}T+>��?\Y	A�>�;��z�������)|���1OO��9]ۮa��c�J��7_���U3�l�;y\~��_����9�v������h���.��xX�/L�:�ս�Q�
�̣�O�ν;Jsf| l��^���jkdM����P��S�u��p }�RR�^��D�`�y�q���FK�Ýv`tH/g�ӕK�V��b���Uw�w��:�zkf��a���G�P�T�oI4Yմ1�2N�ʧsf0�[�Ċ�G�h�j��ҍ	)��[�u#���"t��oӎ'W�����Lzj����*>�ZZ{���6�~���lНK" �2��K�zx���R~��������aKs��ͬN��k�� )�+ƚ�WѽMw�f���ŋ��
rm�7��zf�z��wy�k���o-��z��+lv��n&��3��r���\�L^����������Z�-���L0c�쥶H�Z:��0C=����mRP� b�P{5I��!鳠�0@^�3��4��gvWry��F��	x���M/1�dmrsU�[b��#Y�(�k�1ΦL�p�6]��ؑ�Ѩ�~1�pfZk�A�����<���)]���8����_��h�ū���V@� 4�إ};M�(���Ky�9hv�(�/0v���?4l�k�[�5af���L֬F/@��&]>w����������r[%�9�ĕ� ���_'�"p�bv.������}��+�Nc�f@��>O0����`�dQ�������xs�WŠB�������Efo�1x$rb����+����Jk2�f�H���{��p	���@;�!_uP�i6��J�A�P�O!�#q?�q���q_��j�������;���'�9�W<�.���^�����YZp�/�wL6��I�t�[��1��/&�����Bᥝ�5�O��W�3O�]��?Ш���D~Mo"Y�)�2L��Ǫ�Y�nG�2�JB��
0�[�f0�p�
>8��-���Q6��zg���6>�j���L2~���36�ٌ�E@�٢����_���N;��c
Ѭ1�3���%+�Z���vT�s�Ӓ��q*�D���l� eh�s�j�ʒ#qD��P�4�0�O�z��O'��s����w�ɩpQ���ڄ����
��w����?}B���"��9M���T�m�nW��J�86��U7�ӣfh��"J"Z�T��Ӱ6Av����o7z�'��V�_��6��I��"�XL�q�*]g~�ّay��/C F���=t�"� �O-�|?�N�GlG�7$�u����0���٦OW�/���n�z@��ǥ���W���ψu{*�).*�M�y����C^��k���%��!\�S4P�i¼2B��C�*��m�B
v~��1kχ����[�� �����mF�-�}��n]�� A�!Sl¹
|*\��is�X��5{��)������5�yyn�w���qo�ɬ��	��Lf����`�U�1�ֆ��.�L'��-����H`Ҷ��S}�����5F��L��'H�Z�[�%�߼����YN�>O���=�t�^�>f��?��G�8����_1̩�uCN�o0o�Co��k�u����GZhg��c3��\���M�HU�쮧x�����'B�ƌ;7߉O*��g#�V��S��b(�a�*��%d�d��8B����)Cu���UBs�u�3����~�l������H�##c���.�M%�@p�_���*��.�S[��e8u�����^Zd�B�I��q�]��KvC�V�W��`�x�c٬	����-�l�D��f����1AM3Ɩ�n[�ZL,_��-#ؔ��ry���Ec�غ#���iJ��>i!m�V���n"���	Ή���$!/&aΑ�&I�
Wv�>��s����5B��TO�b����3�ߍ���:y��.V9[�bq6����#��Cd��Ɏ:��*z��N��:�l�-� L�e�{�?㽾Țq^��#��H��,T�|�J�mV@�7"�����8�p,x�u�(�|��ϓ)����=� ˰�k['�ȭI��_�.�C�mFg��S�j������	;���Z�<���{	
��t.I��"��2(�v�8D������I�<=`;���^5�!|��LmO�م9O��9�e 77�6�5��K�BG�[��s{7��`2��\ONz������iZ�<gm�	�-�w����[cEG��l�4�� ����]%*�u^���D4�<�ko�Y�^K��W}x$W�馐�����ݲg]W���3TQr�ɠ�iF�R�����"^I!�Ĕ�wi�~���'�S���Ť�u�����{iDN/�>�VV��d���Hj�Wmd�r��
(J������ͬ��V�T�RI��=��p��d� ��veP�M�|P�����{hRG<�&�`ݜ�}`�
7A=l}}�$��;D��rjU���) �U^w�`��aA�J~CT-/�o+�7�42�����8�n�Uau�r�V��E	P6#��恺9'�v[���С�1�f�x��i��g֍�h���hU�uܿo��f��^��*�3d�={V��d"au�E�� sJ�ekC��-�YfU죶�#�sJ00�+�����Ud�Փ(�t�'J��ʉ�테�͝����t����5rޯ���ihY�Lw���b��r��v���]��X-��#r�E����j@��
�NQGVߣ��_��bGF�Q {qNp��}u��H�[i��>7����bj�H�9�3I�ڈ3d0x<���`ցQS��#����}�����j
+S�-|�F���:�l�Sι��7��V��yi�;��b���O4n��	�]�b�.����4��R��2�b��_���F�kR�܀�:�?������bw��M�$4Ł��nG�u1�x�䞉� ����y	�b�-�E�88����j�����|�@{k:_ОX����256�E��%e���Z�]���B��i���!;�K�����'�Ѹ>$�h�t��ir�2v6l��pQ�Vf���I/�]?��T:�h31QS�){C��(�����%�ȧZ�H��r�焤=	'ԟ��	��>�kL@��ٖ(�EE�)���p�R?E�:���t  E��#oD-�V���8��Bq=^�^b d�?Q�8��	�+�vcv���-v-8�7E��/����e��Mߧ��a��x�
rl
��BR�2moΚ���#\cP�|ޞf<RzA�#I�`�@�#��x��uLj
	A���؀4�P�L^dY����ٱ޿��)F?Ncg����'
ɯ%��������F��[Y�e����&;9g.9�pw�6@�N\.�&��s��p%�@���=#������]�������j��M ���Ej<*Q��o.`��T$���>�닶߶��YY��������DP�ۣ12=D���#M=z�����I\�R��3��V0�M(�9��^ph��΄<�1����Ö`��E��Ǧ�����o)_��f�m�u���w)̓Xg�������>L��%[�+ꩄd;+	�b��҆�a(tw8�@^���q�y�Uݍ�y�Y$>+�Ot��џ�����;Yd�t���zD�ߚj4K�-ˡ@2t'��/t��� ���8�����_�<l���k`��� [�������ܟv忘I�/c
�G&�m���	gh����p����4��/�����V:�y����7��x~�6)��3�j��"7��۬t��t� B�&���=�GBH6�͏�43���}i�*��ēD����v��9�L����ʕ��sW\ L��G8�qmH��"�mc�����䷱�~�,i'o��7��ƈ��Ӛ���n�l���J�fb�?Cj>g�j�'!J��C�+b:%lK D�f�����*3�g��Y��@�j�׆�. ������b��窖گW"����_��Scc�3�%H"�d
90�^*�����S���ڀ;.��9����-OS|q�};,(�m�E��^�V�p�b3._���a��iq���S�[�z�<��9���hl��|�ГGE���0���ƖEE�
��ee�3��􋿐��ƚ�������L�GՍc�$��P�ե.����~���`Ci�i	k�I�J�����{Y�m�V�z$�_ucT0W�Y"/РN·�3��.���7J�E�䠹TF"�^hRA�������h�W���P�X.�*�_6�%�eV��r���a���6rg3�ȆpJ��ThKq����d�S�Tp��9���̥S!�X�2��bn$�`���$�
Pj���i�bl���i�"������j�F�{�]�Q��'�@R�sK�J�d���߽i l����r�նX��>�'?��|e������Y�d2�}�?BzB�Fb ���!��d��'��"�A��H�ա���}��Bizo�'\0�������\@5�9�6�Q)�k�ENQ����e�wy3ɖ��SYn��x�$�^��� �G��d{IT�Y��E�g��馝��T!�Pmj\B�M��fs>m��/'�uE)�ȁ6�¤!��_�{9z��Q/�ʎɞ����S�����$�/�e����g)3}:��I)J�������q������;�)�Eb��D�k��9_J0�1�Q�t��Hq�3@�j�e��j�-E1_�)r��� �-�+�4���؆��k�g��o8[@Sb��\,
[�'N��K�5k�� �G]K�� ��}�%��;RN�K�[�>���/kڂy!��SF��^F��G*��QK��p��_&|�Ai�D�k˘Kq+��hB�RH��X2�/��&n���ӥY���y�)I9A��F�K�L8��J�f���!GI٭��)�&�YQ��R�续��>r�Z$U3d=�x�)�j2�d���;���6T��zA4� �c�������X��(f!�Z�0���������m�2X,��m��+����ڬ;i��!##�T9��B}p�ǒ�l�o�:�7�^"�n��k�WS��K.������(Ψe�8N#1ȼE�G���P��SY`F��sb����NoZ�U��S� r���hÜ�a���:�(^�!�����ؼ2u
䕌״�	�Bp� xG��Q�
�x��]��L�ZQ���n݄���AXS��Q#�J���]+�@��_���O�MK?��ay��q5㊑��ٮ?M-5����ikċ#Li-/r/xC�Zq�u/EJ�˩��$��FȆ��G1AB��V�����/��#e��
�@L�1����ZxKV�X�a�Z���/���xŤٞ����M�r�W�c�C@��zi�y�/O�gPz���E��6վ�5"��hi���HZ*ьW�@�"v^�u��w���Ou�q����W������ �jdi ����������}.S(��ׂb,����'_�:����w���/����Ķ�K��I��̐�a=Ap0}�/�����~�+p �Ps�.���h���=>}���A|2�.���#X5&��� +�D����y�v��R;�(r��&�10+��G�Lc���Aq�H0��"�P���+��C���grۈ�q�Lw�t4���@�YK���LXv��`�Z\�k�s�b�Gs�Y_}�N�-,�Ǩ��I5�'���E;(vÚ��Bn�u��Ӷ�'�i�8�}��xj-MC{𕮠M�`p��:6X}t��r%��#<�RoN�m��"J�xz_�(��!:�ĽXRH����ŷ�Y;��J��6�Xؓ��.\*����Hۢ!H�	{�F�'r0�X��"Z�Ƃ�6Ͳ V*�@�G�a@�"KcR��!��z������3����:��\rwe�.vf�ݭ����k�uR/���%o5I�;��w�,Sx��rv��k@�&}��8��� 
�� S��D��Q3G���R�P�1:�6�QI�$j���B�/d�]�>���8����b>��a��ErWO���Gb}u�eHȤ<�-���὾��4�8�z�����r��n� O�bmIl<�uj�X�QZ��3���|��ԃ�[����+6t[ZTM�v�3�(@����Gn���X�{���h����Jss�@Dh� ���#��?,��'o�HV&Ǩ	��+��9�D�RBSt�>@�����#5�\�B� �b�+�1�����AG�'��2x%�w8�'�z0鄁�d�O�����&�Ug?.���7	$g�����&��R+Wփa�_ꡮpi(��F�W��s�%,���ʸLz/�+�ܴ�{7��>y�1oWx<�v��J^�~Z�S(9f<�~�b$�o���/���� �)~H9�xU�:����t��2��
�̞^������ו�Kn%�u6p��1#��"�.�*�����*E+�D�~�B�#�`�o�Z⨃0~�R1T?_��uBx=��6�0��+d9|ÍP.�6�ynpq!�|g9�
��D%���fJ�B�'��dލB��9�J�H��Ce�8�`�!�4�ER]��VA4B�>{��r�H�JJ�Q�+iuid��[2��֕���%� ��.�gY����:1�I]�Η�G�D����$�B��	��	K�!�h�\��g�fZ.�gr��]K$3��+�y'��ݨ~��ʮ��n��6I���cB�?wX��o��� �j.Ӧ-�Y_�G,yx�@�8�᷶^�%^i�����fhE�e8�ܧ��Sh��c5q�+6�H�̎�0�L�s<?ͫ6�r�W�DP#bN=��N=�ǵ��E0�JWv��y& F�r�Y����;nQ!M��"";d�� ��Q��2�DץV�Z����͊p'�%��(���KH�*8�k��;�Hn9l��hӹv��*`Vxo}qݏ����c���"�)�v����Sw�7��łux)6�T��{T����{���.b΋��b���0ь;��t5�ئ�z�xH���LI7Z���@,��DF┞1s��Ϛ����t>"/_R��M2����)���g��ہ�SZզ\z�I��=��6׷�|C<k�d*�+��5��`�D�tM*�|W���.Di�>Uk(P�	��n �:���'8@��,S}�6pmĂ�>�hW����i]��1�(n������1������[[���8�Uw�"�	�[YSu�;.��'�,�Z=[�L;�� �������*,��4�7��h�W�H���� �r���(�t���i�"�ы��$=G�ʱm�vb��S�Y�}>2�|���ף�^��q<Q� ��˥�G|/�����M�NV�^yN����@ѷ�]�����N�W����Z�ؤ�x^�_���D9q�a��n���F�GY���¶v����������m~�g�R�Չ��;f��p��d��,��H���-�[uǴ��-[ϪJ�*!��Ѕ��K9���
QPp��R�s�'�H���CC�������&�2�m]���|:��W�,�Lϕ}�����q&�F.��U�ږ'�>�i؏k�[�!s��f�rl?R�ږpAƙ���\*.�˹91����]\��P���{v�Z�ar�Q��]�%�V��dޗ^[��"%� ����p�6c��E��T�8~?|(��M��p/����� }8N�#�Ji	ұ��弁|�ֺP*t��Ƴ�v߆��x������W�OjC2���;���{��+��k�l>H���z�LG�D�z�v��	#�j/�A�x"��
��k�Sɮ�>YcN_�ۥt/�w��[�%�6�m�����I���F^..����v�Z
�����A�k��S�.�e_v�5���m�!��_�!�=iS\�7����j��$(y���u�p�A@�7�3���D"}<^u��[�oł̿<��k@,ӿEz�JeBO��;s�+&�*��f�W�M}���Yx]����,��o�Vtm Un��o/�k��:�������������֝�W;'�Jc�F�M>�i�Td^9}�7g"6�-�$�s���O���_��y}��M��s��!]Z1DJP��PI�B~��2%�@p���*c5�R�C!l���^���}��H�jfb&Kww�]����������C3TԻ��H}���O�۴5.�X8a�D����[L�u��騫�l֘�C��������:qt:�>:�^��Q�yb�<�n�9�	��t��|G���������,}G#��Vh[�][��j�I���q�PZ=�:����]ˆW�f���;$n� 졐ײ H���Y�y�SK|�Е:�$��Z���.�o�^����Z?}��ް���eZA�J�e��G�m1�y}�[���?�<����c�O�E1�Wņ��j����s	�䝆d�C�����&̝,#K���~c��30�gZ���L���~H���w�}*��?ʆxG�hgK�C�ܨp�D�� �t��.+������ǅB�r�~huǮ�O�@��զ�F*���I8X���	eG-a?��1��2Vt�t����r��� ~��\D��N��)ҫ<|x�BW �n��١�iְ	� x�����Kh�����-6�8�m۔o&�������0[/����B�e'���o�<���I.cϣ����*l�T=zL��������=f��StE��h���k�j�AA�8�zL1{��c[� G�|	��>�ځv8�~�܉��d�2����7@��R�3���3�`%�p��34����/r���9����@��^<[Le&*y�+�h�{��[��ׯ��#AY�Dh�]%��t�HF'�SK)p߸�
�� wmVo�q��&k=�Jj^X�*Ǿ^��}�].��h:�S�u���kL����qvg��{d䵘o���:.��D���5Yâ?O� �\qg�Н��!��,o SD?`Ǘ�7�>	��`�M�������  �3�ʳ픓�R��{\�#G���y��x�듚#��8_�|���K�*����d�ܬ���x�!q�b�g���{=�w�L��o������10����h����Yk��,���q���w}��O��P{Jꡆ��u5�-�it���3�@�_8NeE*�E�9ސ�3u?�W�X��*���cE�A��R]D��>dV-}:�p��?EIGGG~6,	�Y�R�/k�O��ȽEk	H6?]��p���:�Ū&=��E�;�A�B�Q�zL
�H��. �ָ�I �SXLf(�nW{ ������ͽH*�rm\����Y����_:k��rD�Z J�Ψ��F��Ԫyڵ����axU��z�>8�L���O�d��B�h��E����7�^�Ň�ٓ�ڞ���AΞVA��{,|28/%�o_�'M<:��[�aLZ�CM9����L>g۰f�\+��}r%^c�K��ı�kI[��N���'��<�?X�B���(ԉ��nO��Z�����B4,z
n�_�����u�&��>��o�H�-tt2��vڌC�ç_2���q/N�|�\X�hZ�!@����0/Ņ.��P����_;SX�0�$Ib$���LC���a�f�0���C/�-{�yW����M�*S!�?ũ�~E�|��o�" bż��w`�:�$�vx��~�F�
j��="h����u����4���Դa�]�i��7�:��j�A�Y?=��9�,��,��Pە�r�:�K�,��Wx�����Ag��D/�=���~d\�h�$�LEѓ���5��jG�g�0$(��-�������Mj�a����>B����+�P-E�x�����7����ѥ��/�g�g��˷ɅkI���^���#l��׈��t]\b�3��ѕM*�tFw�����w�1�Q|�I��"8ג�9'Zb�3�\�=���n�Q��~�dCs�g֕p9����G�qf�5�Bz��Ƽ��]���G�	A@�O�+�N� �1&)\��HG������2!��-���=D�o��k�h7/��������$Q���M)E�ҁ�~4N�c1x���{�$˻�`��GvJ�{�XF�`�<�m�� wT�TG��Y7�y���׵KC������������(���Dc��1)vbQ�iͨ��
�+~��A*�{��/I��f�G���O�/_�Eْ�����r�PNs]�w�~�Ǝ�a<BЕo��D��=�p߽�Y��P~��K�S�;��~�8:uH5a��9klu��[B%�R3C��I��
���d��I�՚�ք���VV� ❱љ��G�����7>a҇g��bcR�����0�b�ӥ.aR���Akz~�Y1Sw�q�� �91+�sƩ�A�:ůN:�N�zn�	w�P��-�=?����ɇ�Ek$�S�HQ;�y�Jp���h%����ۼ�`HGb]`
�T%������o�fՓt�`/%�)c�}�#�i ����'X\�*��X��h؂���3�����N3D>���7bz�y&�6�6�N��9���S�Kq���0�#J�֌����7�t��XMrqB��K����~ �jh�p�3�]��M�Qyʃ�5����;�Υl�]~~�*�B�Գ �yp������bLA�*�;��"L�}��\}����E3.}r����&�u��)�TCG?X�����v�K�$�/{%?��~�� �XÑ��44}~1�ÏlA�����RoCG1�� $vC��[vbf��R�uC����<2%Y5g�Uv�K͜}��s�,s��z�80yx�"\Rݬku�zC��!�\��}X���t�ts_4(�uP(�N�'}b�-��OXU5&����(�u������lo'�i�GE֣
�4mw5l�R�ӓСq_����]x�S@UkQ���n>ʊ'+��J�D�}����	��2ϣ��=܌P3��Vs���������m�x "w`l�#�>̏�CW8�C.�-:�%E
��%λ�#�/A5x%sQ�*�� ��Sp�.�]10{"�P5ǋN?Z|���TT�=�/�Q����i��8>>�!���P<a�a���h3�����K��@
=;G莉O�ud5�E��y�	XЌ� ��`T_�7M�o�D�R�x�Zf��	���o�g�A�7a� y�S�6V�\��0$���H�Y��$Q�9ښEĒ]�|m�����)�F:�\��D�Wۿ�F����	~��
n�W���Ru)�@i~��K@�[�˭���P�%M�r8��|b�u&C'z �p�5h`	[y	��S�Ԝ��������w�>��=$��-	uU���4�`�֘4�i)�L�kS+,\x���:4��總��2]��@�)��B��ܼ�P�У޶֞u�r�4:��'�ԯ�Rh+�2w,b�2	�yeXwo�3�nl�L0�ZW���y��i�T6�	c�ҩ�kAyQy��6�'�EI��c�	`X:!�7����R�O@�$4-�x�t�
}�Onƈ6��y��H�����mE�	��W�N'��xb��j�T�p�f���S���E5���w��8�R�0��������~x��[Va�_�.�G�ѓ�7���	��%(%����Ac���@ۧ�g��y����� �Y��S�*�\����!�1y^��h�OT���&�RN��`���'`�o�������?{�ZX����M�l�q��������7�sZ��}r�jTx"s񪈻O^=A� ��:�J��lI*#@T�+:#�ݻ|�>�xo�J@�2"�[lq��D�͑Q�%Re�e4��i����I���|*�hY�5I�����9[����#�����w���6�b����U2��K�Z�o�I�H���m��S���.I3�K�d�NFb�9U0�n�?�<8��B�;"�V5&=I���Z�Z�e �N&��?7�d�9�Y=d�q���]`J@wھE����5f�&�d�Mus@�0(�|X	/^�Ph�5Bؐ���CF
�:�z1��&��o�ן���xGA a����o��}�����y�׵�,�αq'ޚ�HIBҧ��ZYT�_F���>��Z��9i�p[DT0�8y/��Gq�>�_f��M��*����/���`vb�<������鴇s/�}�T��p��#��u���(�*;W,pv�;��-l$���+���i�\�'����EZ���~����ځ�Yɺ��b�]�]����WQtZ���`��
>	\NC�=�����&����X4ׇX�mn>vĬ���P�pяM�.�@�b����*z�-"��5@p��׵�+$��yҮ�0Dz�{�v<��٩�ťO��	ZV�m<�
���tҚ����&�?W������>�R���J�4F�Z��C�=z<~s�N.vy}�C��gq B�8��uª���� jJg�����荍s���u���)5��E�C�_�"u8F��E�x��ԯO�������,2m4�O�v�f�a~�EjWMG�"�xF�P3�tR�(b��s"��Q,�t���A6X���N@m�p6�!��
A��<� $ n��gA�?p%�&�9).��9!��P���O�f�?=@��}Er.���D����w�6-�����},���"޸�nk�m}�2�.ؙ!b�f��_яF����Q}&��֜�!�{�ӆ�TkHS\� �(�Ik/�KK_�Q����~
{�ݺpt5j�jK#��]X&Ox*1�.�&W>���./�gj��dK�ɱ�L�V��R�	��S8�j3F�>�&U�	K��n�~�T�Y ���j7��'0�͹�V�S�����=����*	K����]�s#��Ư�vA���m��H"��䙾�_pk�����YƯ`[�A(��H1�����ŏ���<g�	�
��R�N.�%�<G�[��u�`,�%_^ct'�jtݍ�a��L���-hI�����a�R;�
�����N�k���X��S.�`B.R�d~��nj�m�4	�2��w�������1�^8a*�u'D��~7H�����#A_�43aJ^9���2�������@*���0\�������� ��"}1��Z��A���FO��(7*���m��Tq�N�H����X���
� Ȩ���h�jѮY>�չ*�/^���_T��ը�D��ѯ�w��7����͏�&��#t����C���b����r��+�>¸���[����N��������>z?1��L�uO|QҖ|�$��J�o�RtP��N�^��0��2��+�b�~��C�?���ލԻ�R�̝m�rb٥�j2Z��1}�o�A�I�y������ԋ���}�t�~�Ĺ�Ey����uL,��۞�Ŕ���:�Сh9zI��g��I�+����/�>�Nb�G�g�0�-��p
f�U%�א�i)]<�Q(0����A�n�F�U���#���`6[��|��wr1��(�������b�?w~�^ �Д'"od�a�D� �H�TY�s]�X�.N�<i��4�?eJ����ϊ�� �qFPU�XO(���3$��k���DKb7r�|�
���8i&��`���y���,���-͑Lǥ)>I��l�C��t#:Ӵ��rl4��?"�fEh�\��E����̿" 0�F�B�)A�����肌�x��v���\�pI���ZU{DU)6�&�<̈́j1��5�2=<��^E���RV��>��9�\�3�yDqgD~ş��@tB��׊9v�Y��Iw���m���� �,������zx�?w=^��4�:;����Wtʘ�����v �
:������έ�r����G�z����[~zj��� i.-�[�5�����2������v%wNx����6Y�4�7o����8jj�T��Xކ���*N�}A�XM��	5L�(s�1�d��j�|IY�]٧8�&�L߂؄���c�F�cO��@v̤��ep��f���{Ѷz7I����N~��!{I��B�Tio�u�o�'�/Ur�NJ��H`隴@�0g�_~�q���P�X2��y=EU+�Jb�R�XO���#C�������x��|�=�u0^޿�F��;��\<]*��ͱ�י�I��H�l��JT�4�(gd��q,��H�fr(�5���~���降S��Q�C{����[F�	<��=K]�3{@ b�tkdy���\Y�NDȘD�W�q,Q�[�^�����L����N�c��#U���ɰ;q�
1�1�jYtx�չ�Ҳ��j\�.[̞��9�|hG!D��%/f"�{� 7�ٗ,t�(x咘/�`b���1���|��@��t!���ӦYZ��A�wS���|��\ A�àn+���b
t7b/AX���a�Nͬ�,_G�1q��z<s�����b�"I��������q^�x&��Y8m���a��T/Ծ�:A*H �F��>V�;�n�[��j���'ҡ�������b�~$q�k�����᩶d�/V@0}n�ͬ��6.�lnb�J�Ze#�!/,�~�Bd5����;��$r�ǳ�:��� �ݫ����#W;��'�S:&�~� 4>5��h�:����k�*"3eR��g����%_w57&����&�{I87k�����X��f�A�ed2ѴU�9p�s�3Xd]����qڀ�ikW(T-;�P����й��LKuo$}dN�2�e`0� z�щ��	Zˆ��AF�ٗvt6�	���w�����`�k<�����d�:k����}����l�1<�va�lgT��KL��
r�O��z�F^C6Ae�]�32�C(?Uf�^�zA�|՟��~cnn��dT@������2z���k�4L������{8��@����;��~s&I���v�Z�9���ar�̘@'�aZc Y�{�ӼU����wZ(F��p��@]C�6��*���l���0Ү�^,o�F�!U�.R.+�溉�%��*G�%�J���*�u�L4��_0ec�8�P���%"$��r�����;!���"�2�AjBpʩ��b�띰��Xxa��^��P�{Q��"���8�	�ї�{U�Sƹi�8Ib�h���%���#��7�֟��GЅ�3���@�]�@�ͫ*|ç��]�V�'��m��FQHR&d@�d�q���<���;TaA�g�skqPw�/��|�(2v"������=�������u{?.�yLĳ8��T8�-Q"��&<C�GÒ{PL!�^����3���fW|̎,�B�!��s]<���M�<�m�陎�HR��~�w7��0d����Z�0�P�R�.��?w��I�b�9�br�PM�(�L�Y�s���(���P��	!��vP�KyA�#��B��/=u�����`�����a������^��YN|��r�(�pךS���n#�n�l9�<�n"�Җ#X��G0��*�5>wXV��:��o�mv��;��}�-���H�B�Z���vdn�y�^ӧү��fw�5������W:�g#�7I�e8p�A!j?	#p66�,���k�EUu$�Ux�f9u���č�u�%Rz��-f\�u0���3�p=�H4�����l)�e�6����p�ܖl�Ó���{��������{;b�5���(uP�����@�c�yx�ۢ����"�i1�}쪸��2�`�N�?��"�+}�_1������xx�4���b�;Tq�P���k`39>9+�}�����i5�ή{6�_h-����r	����ᄄ�hK��e��8�_6ҥtex�d8�GhB��@ɇurl^���CRK��I~PI�id��)&"����[�*�G
~�ƨ�x���)%1*��W���w' ��U�rV6~���P�z-����f�� �i7<	�D����
w��D�����ц��lo�d�b7����G��mgs6�]�oO��5쁓e�����J|3������ϊ��(jނh� 5���EO�-V��+�f�����Vc[1����+�6-
zw���D<�R�8H؃A3��v_\�v�l3�T��/Č�J8{��s~dR�(+�y^�_rc�@^Н5���Cݝ"!J����Ō-����;ᵜ��2�A���0�<X|�����sP ԗOT�k��V���UD-�IK���>�Ӻ����"��q��?w�UV��uQM�P�㯐���p�f9h��m��g�x�/�c�œ��kJ��u�*�|�(��G������zx)]����l��3�G�`bBO�		׽�#�jLU̙C��1�R��U�r��̵"�W���q�
^I���cg3$D��{]�=�����hى��-O�d�j�~ �d������?�A�Y]����Ԝ�J�&Tp��t��p]s�F�ES����!>J�O��/��5��F�$>�<��V�.�
�)wUoFn�ln��<�6��0PP�H�����%=���.ؚ�\���%q*I!3��LN<T�Q˰	j��EǙ�(?#����[�����*�X̺l����z�}8�T��)0�B�j��=�zb�<*����MmR!'t�{����qF���1���`!c1L=ݗ�_r ��N��)��`|w}�$�/�ǃ���U�[(�K4��`x\��LY�_o�C^��2C�����`��������JB������{��ϳ�9sTD�=ď
:<�o�nM.*�:�!�*4{��Y�4�l/�q���p���+���
���L��ک򰲆P����,�D���ϟJ�9��$cz!��M��Q��VAvZS}�^>��ßsY��gg�y/����[c�Ӆ���N+���{�6�����T/�'��oI���,9'Ȓx�B��(#u�v8"Ž�<��s'?82�/<Ip 1����,�
�C��,AH∬"��'q��à��6M��v�?�r�ݷ�K�~�0����s��d��ҟ���k�c���Bg�<!C��3te.dj7߆�Zѡ+��y�����M>��B�|���G�[�0׸�`) �����/L���0�W�:�g�x�C�>3ne^�
�j���:c��D!���>zR|�/C�8y�.��N*y,7��0�S���uL��٨�7�_�l����������M֑����Dn{4t� Av�ʆ��8 華C�h~�H��#�/�����r�Ы������:�I��h��|�k�����I`L�S�*�P$}� �qy��i�u�j�4f�(��zlN)<g���F�O�`❧��%UQ�����j������J�x�	y�?r��pΈ��|}k4mX��&�F7�@s�ݙK��_��x��,8��:�P�|FG�t�����%`<9��cj�tğ23	����^�ȓ��w-�8��kωBH�f�JL.`���a�x�LM�r[(��Јގ�_��۽�1��r�؄���vS :��e'C\]�B����g�����f[Y�XiA8���*3 s�b>�	�Im�v�B�#.wМ"#5NΩ��B���Bp�k��c�	��fcp8Mޫ|��#����"N���;�Z��x؉X�{=V�$K��������׆�U�l��Ř7|�?Ƀr���A��3����א�ڝ �iS�A�Ɏ�UM�ò�W�h2�_�1����.����Ɓ���!
�c9HC�����Y�����]ΙL(l�c���X�H�<�A��x���,���4����a��%��)�rܛ�{�%a��i�vj\	��R�h���6F��JJ޺K�y��W��$A��J�ծI��U�cV�����(�A˃՗�:l�P֖(Ma�,���KJ��+��{���鏋H��Wm o�:u�/�t��ڠ\4�;q��jbx�f1=KĢӄ����*ytE����c�Rb��"�Q<
�Ϩ��j�\��{0��`eS��W�I3^�C��G�io\����