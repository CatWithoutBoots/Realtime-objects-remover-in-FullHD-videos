��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&r�F���oh��m(�ʉX'?����E��fNom�K����[Ś\�������tT~3�OTA����֙�s�͔I�%�@Bo��H:D�ޯ19R<h��IZ_�?By���^X����$Icu��5^ܴ~�"�=Li�¬`Y��i�X�r�G���0��*@f��̙��n�ʠ�?���}�	������m�,
����
:?+��J��C�4����_v$�f��R�,�� ���PN�TҔ��A�*mxz/���Eu<�GR�"�@�]O�
ǩ���ļ:�PAT��آ��+�c)��U�%��E�D-���#Xp�(��P􏃊ñ��p)�@��W0�3�Z ؐ͒d���Q,:��N��1�+S p��e��?|N��j�O"̯��pp%��C�q�lō���x����4&�+j*aʅv�09�u���D�2[O
�i��D� Dzv2�j����0�Y��������E:G�����4hlH����Z��Y�ሻ>�D�zn�d�B�|;�'��L��<g�G��K�?�0Nz^|a^��!sXn�8P�m{q̖��� ��{��֟�9�)�N�����_L)�Wz�}2�L��%����=�H�tȴ��[jU�E�k�&8��,�/�u�SO���O�$g�lZpG��R�I����K��2�pD�J�o3�KNj�w��W���:Ϛa�l�{T���0�2�k���`��Ǘ_5,5�įG��2�)H�W���J5��8� +��	���>�X����'J��C���~���6-����{,=D}����¹��B&y#��Y}^BbI�4YRB&�?�h� Ķ]�`9��������c�E��/��E΋��/G��������%���La7Kk�Oy0ߥ>̒/�w	\�r��(Z��tÒ�n��V�;�ߩ\�fb��޶s<<(�O�X�߿�e�}���x"�6KI��'nV�ąi �<�O�=B2��Iݸ��аr�wn��(�&�'e���eQ!5���=FtM�����-*
�cǿ�qm|8�ަ��9e�1�I�[�>�݄x�f����N�!�C?fC�����jݥ>cgZ�ۨM,��]abX��vRy�c
^��R(����� �����n}F#ȑ~+:)�;(5 =!0z7#{���w���׀w�d�f5�ͯ�ۋcD�A��q�H�ś������29������
�W��2|�?�kp��ƃ~R�#��]�gJ�Z!b��n)U���g+_�^n��V��!���	�o��bӀB�לkD,���Q��oW<2�����QY�+O��sH��A����*��cO��p�XT���	i�� ��u��Sw,��8=?����X�*>K�ﲙDp���3(9׼��b�3�78�J�rsy��l�J4���m�M��%S�G�{��[jT��v�����;�@���S	��� �!jh�t+U/3薗�K�~1X���T��)�_Qُ-Iu����9ˤpc� v��3Q=@��4ղl�X�5/.�R��7�s2�5���is�u(6i����&�A�k,M���ҋ��RN�!I����aVq�E���H��X�lh�=G����A�:+
�n؀�s����P6u\.���C��\�׬��a���`�]���`/�k��c4sΣ$���SL�*����Bb�쿴�;u��wf&�:�9u8��}�nb�NQ<r�L�d���;������-�'hF](��5_4ރ;)�+��6+�2*a�p|�gn�GP�
O��(��(����9�{�N�[2x�M���lZ�?���?�c�F���r!���u���IZ^����"�/8K}:��A�>�S��!�R���Ap�� U�eX��d�7��a�+�PY�
�2�R��7W*��-�%c��Q�'�����>��	��r6 ����!����i� �F�q��3f=0��L�)�c	�(�j<�Vk�ɶ��w}5�l`��<�������p*��PjԃD{��(�3�%���2�zEJ0�0ɞڽM���I��S�p=��""q�(�ڞ��r˹/�?��#�Ӏem�I�@�P���B��J\�ok�r9���!�����LD�Qo
qZ��1˯T��& �^��d�86�y/(��ëKZ%�e��,LB ��!�_�6��K�83փ�DeH7���;�3��-@���}N�B��ZHҨL\Έ��J�f�x2����0��Z�/UG<��Wn�� ͇�[����!���xP��	.�[�s���n}-cTn�?��\4v����r�O�z�X�9^�v.�`\��2Ǌ��0�Cnγ�?�v��=���\�R3�Ppa�����9��������s�i�6/5���I#��RC��q�o��
je��{EȚ�^lɄf����� �RG�S����`L�
Ug����&���0�n���F6ҟ&���S��E�vŐIi��u��gZ@9��W�V 	�t�d���d�����q	�k�XB�Hu?/���܍��w�)!,�\u���+����}z}��P;n���C�6}0�O���6wmy؋O�pMYa����<�U�ߦ�����»9Dj-Z"s�(V3��A�c7�)�ů��_��/4)�f�?��B�>�(��!w1�#j���J�z�X�d(0�ym������Ɇ��Vcm�:� �J�;�jC�?��q�K�o7X�����]h���z���r�u� �Ҵ�͟�=�
R8��rgi3!_䅈��<% ��1ٌ�b�޸Q�4h{�\��W�B~����67�Vއ�a��h��ȘǕA
nE��'�F �B�P�g+b�S�J�á�0l�@�Dz"�O��]�9ν�MD峣��g{p���D�	/{�, ��\0Q�:�ɠ����Xɱ|wZ����,7I�foE��J^rA�/0~����LƑ���K���B�4��~sQMT'�<�v�H�G1xC^i��|
���CCG`�vy��tf�̍��|o�{�=ny.��!���!.�3ic"���,�U�~��� G��e\���k�x�#��W�hh�	������p����!�U�+��^�Y���V���/~��W���؎���,���7�U~Φ/��R�ˉLC:���c�M�KW!>�����Q��'V��"^=�ޖ����|�.��3h�7�g�@s'�A'h�o�bx�iI_�Z�o<ĉ9�[g��s�7l�!�'D�M��"�c��B���r�r����*��*8֍ڔ����r^`����a2������;F*���Ӂ���K��n��v�� X��?t�x�p�j1���'�u_�h�;E: ��w�
5xW~Q�ֵ��ϸ\�詐�������L�]��{�k�"c�weon�FQ�����u�3u���H�wW*��ID����D�(F���p<H�R	��e�e����^�{Bt��Ut�_UA�q�@P�I��Z��=~�^�9Q��6��,%��| ����x�s/�o}�t�V�!HM��M����wB�s$=]�� (�G2X|��6b���`?/Mt�]�t{[_�]��Ø�{�3���S���W�h�_^_���ː�H�C����|���o�v.�<|�k1m��ld4v��v��p�e���j����A�� vs!�B����9�x�W�����	e��\_�fs5pTl
p��v�).ܹ*��j�"٤�XV"�$��B�X����1:�U�c �b��F)V�Ψ\�e�����
z�'��;z�9W�J�@���"��ֵ[MW�~����rT��1߻�	A2U�Ԛc#Q���x,�F�x5åz}�cB��e����j��#{O����*�-���m��_c�L7ͩy7ō51��r�[��^m`c�������*]g���0��nSG��ib�[u�.L��0�#����7�dUrG�m�h�ܤ����&:N��S���VU�~�fM��`��4ѕv�C|^1�p�Ln ����I�ކ����V:ZX��엷�lHf�UáA�bkZ��B �34�����C$�
t/3|�J)rA�W��+^��p�-b��;�)��gQL�9?́�'�>��T>�o@�E".J�����z���+����w���>�F:��}��]y�8�������(3��+jm������;7��i6��1��-qtQ���:#��nk�v`(�7H�s�g����tϦ$��Qʓ��n �T~�G��^a���R��8��Ļ�Pgg�-�琯�R_��>^AB �iU(vQ��3(㵠 ���ǁ�D�kn���@���M��tU߲�	�!1��"��ة>��	$nJ\�U�{ǯQ}�uj�8��@��duQ�	����]�w?B��\i��Ky�����RbS�@w�{'��
M�-�m�� ?F]I�}�r8��\����p�.�+��D/a��C-���J4��
�~"���lZ��K[������sV����"�eg7��զ�oK��[*d.$�0�<����&t�T<��3F������QǮCC�=-0���W�\\�����>��.�+{~�C<����m3IzĊ5 9<-��o�0��������U"2��`H�_������'�o2����z��жi��E��I"B�o�v�B�����5c)��W�W���d�=�`qշ��ǿ5�U�H�٤��M�/�y�%�._Kg��#�q�P놤�fޥ�:�I,�Lr�f�A(af㚇�ΜFK��#����<$65�]\F�u���RfC���9U� G۲Y��gb�.�kO,����n%�\��?0.��	GR&d��H�zG9o.�<����2a�:���2�-{>2�9�P,n��#VϲAa�@���f��W=���,�EyS�MS�?pآPF�9$J�t?�WN���5�8w������ {�*���ᨧ��rΚ��v!����A�ɖ�}٧���S��9k�r�Yw��wl��a��j(���~�?�B���@[�kPМ������
��W�2�	l�g+^��{n��i�˙��l8M���R��+1A�O�#C�UF 6C[r.���ʨWB�<!�Z�X�GW*�L�9��K�_y5n-Km_`��>H,��`7���U��[�{6ߚ-jN`��1��ayf.v�?3������L۽�(G�@S�>R��S��\�;�>q�4�:�(��DbVN.�6�A��C� �;�̭��9D��D���Q6�1����ދ`�U��A鴫Ϙ�7��j����w�	�:���P�w�(|x�e�A�U� ��^$���B�/.6��t{� �o��Eq�Oε�����PK7o�O�#o��}es��͸�!�_�����Eb�^��p�*��(����E���>�6�X�6�g�s|㍵���QM��1�%�������|�j�$\5>�Z�:c��{r�N��?Q\?�5��O�HO|�1⮘�!Xxn'���Y�&ҪqV� �-�O"����L�vg:*q7u��GG�S���!����)�vo�m���>�Ү�ʑɻ0�N.�=�_ܛ��3!����ɐ��'�*�m+T�7d��´/�;�&b�mꅦ�|�`
�������r&������\5X\��Y���r+|&��=���������`�g���R� �1ۅs���i(�ۍ��
�G�y�ݓ�@�1jDJ�eh51'*?��� �Y>���Z(jo�������d
=S�Aѓ8��w��L2H��P��!�_��i��<pX�����I7��C=�wi�n��CCW��@�ۛ�ϟ8����R�>�vO;�Sδ���Ѭ�垭��Ą<÷�i��v����d&o��Կ�������%Zc�U�cBN��I�z�kMqQ!�����) �f�����nXb_�\-��]�8��9:�z%�$ZI�>s$r��i�(#S.6��KJy����q�.���z��[���Y���S�k��=�h�9�Z/��[�a}����M��g��'�mKp�����Q��uʐ�17���n	h����Ć���/Z��Ȼ��▪q��ޫ~�R�3N&:�ՙ����-�%�RciԵ0i��g��A%Q�����9�{�Nz�=?A�e�NM�{+�6���V��J~�I��+ >hG��Ǯ�rwe$��C乮�������d�@�xa�⥘h-����s(���Nf�D�"�.Ҭc���%|/�;�������e3)D�_���t��	aC�4��Fɴrs��<^���L�\��VUg^���&�JѴ�Eϩ����Y=Ϋ����Jjsj΋>�Z{�$��2(|����6D��v�5��C�<T������i��`W����Z[1$��ȣ�wSaү+lk׳�k�H�!�1�� ��aC#>ܞC�8�ƥ�D���*xhp��e�������]����3	>�!�/����e������v�)zkcu������s�a̾�$m�!�^��Drjlء͖6���7|�9Nr��l�� �%��_�9���3���]8���j�pJ�a],3jKWٕ�U�W�ӊ��jn��U�[��o��*ͩ�h�D�+�8���j�l%��u�I��ѫ9�쟒��{ ΀���ma�s:���/�o࿄r�Q�]���v����(�1�B��R�%4��&�����#�D�p�!Z��@��~]1|a@��I�MH��`�0f��QE(�mIϔُd��O��������{P����'��v�M�$L�_�����7R	J\�hԛI£��ܙV�c�k#P No��y�e���{�R��dB�����/�@���x��/�N`֘��<�ԗ���fo ǳ��;��Q
��g��!�uq_�[�x�%���?AYz�~��=�v�U�v�}�ׁ2V�)r��J���� ?�����U(�A¸���U�e��R%�Sq5��{���Ń���K& w����')���?ɇ}� �Z� i�����M�-7��"=K�
A������G�s�p��r�Cבs��A{1���o(#Q/9&M��r�+�yLU��CjQ���ˁU�����b2:�r�,_Jbv��kC�}_��ւ����W�n�H@�.f3z�d=���8�`L�J+�[�m���hyCR>�8/��
p+ל�%tDE��Ux"����a��q&��B�uZF|�-���D��UvAd���
�u�	�Ij�1;���{5M2�C�B���P�<K������o�0���`͑7��Hf5���^�N�l��?�M\T��A.��F�z����X�Uze<�Cf���9��^[a���A�FP���ŬƗf�U�I%�3�=m�J)b���L�1��4�a���vz��/XǼn�m-�*s��k��>���>�M��`�Q-����+�;��Ldֲ>�����ܛ�k�[�A<��}�����|�1Q)���g@Æ��眷�l�7{?ÓJO��#q6Z��f�ho�v>���Y~��ew�f�uG���VrT�����S�P�c�}�ޫ��+fT��F��`�#�g
"j3���[����zDոc��i����in��f�=���y�Y���`CL��\����9Z��\�-�S7�M�����7�;��8Aau�๣�ʱS&�j���c���ti�t�C>l�I���-T��܀�B�#WP�V,%ctR��f6���N�`���Wň�2JJ=�W�W�Z�+�Y��)Z�Ե?�d�QQ��i�瞕�?�e�i�q�t�ν+*#�g�/�@<>�3B�����>����<=�!�2g��Y��B��h�;@��Ղ�+����g�(�kL�K�,
�[՟}��K����߷?�i�%]wK/��F12���W�vG+	+� �<�j�I�k����	OYԾ����)���Ôk"!w�|�]��������b�&���Bb��r�]�25+�Ц�$�4��=�H"�'�s�{\�u9� ;޳�U��������R,Z�t�LfF��k�C�e��g�{>[����<=#6����u�~��\&B8��[o��N�e�+i���aY��|y?�-���W�E_�@n=��xp����@Fg�9����><�T�c/��s�W�CU\�@_킔�6۴i���p#���g+j~P�z|�-o��22?Q�;A@"���W��z��Rf5N&��۹B��fD��UP'�Oa�8��'(���:�&���hTI�I`��ZY��g�E�g�*^�qQodD\<�p����B!�	2/�Ajk|-��i�Kz Z�\����P�N���q��$(����8.�:�F��:��#����p��s�2�;ݬn��<�,4�$V�VFm����7 G��<����2�p�|�4�c-[n'5�)��W���Ό���{?�ԉ��L�@c>��݅�)O�4��Z�x�FGNfy�ꙏU�U;VV5�0�,$V�s��A�1������g������e!�Q?���9��_Ww���@�Q�����M0f��䦼��h��6o�d��R]��6MU*��<�\oU�#���N����qR�)Xaµʺ�
+E�6��$Q�Yt3�m	�e�����s4_�jW�-k���ڈ��| *������JJ*�����F���|�Tȼ�1��6�{�P6��K*��,�jF� �p�v~��S�&%��0 �
�z������YnǒL��'v{�b8��w�����mO�	�,Wi�W����ɂ�;J�O�ih<�zE��a�6:��͇�TF����-X�8G�)��W�Pi6Z�w�=�B�(̧,��L�F՜4���3215-%lxܳ�]�Mx��6�^�pր���B�X�e3Z��\+���N߉����8�����ay/�^A����s
��D�(��z�?r�)UeF�H'3��_�`�B�޴��$e��X�ovi'�$�PD�*��lM� �>7Ŕ+u��_&s<U�R7���)%��(�p���/��C�gI��b���̏)�K�o.u3�d�e�	�Gx���Q�qd:�����d�]���t.� �_�W�Ό�D�;��Ū��֨#�Hk��ķ���q_� p�l��ciW$��*�~��{���n�c��{�W|/�PC}黇P`9	"�r,�Go�l� �I�<�5�x���f�%��IC�� L݌w���Z�J;�i�˚����f:��B���a��ٞ����l�z�l�:iV�J���ދ��0��8���7"�N:�����w9�ǋG(��5�h��TG�1�Ol��-���J��)�U5�S�k��7�Zf%�vui8ޭ1�9���m��?b�7(sS/7��/�{O��O��3hoE�%^���F_P}B��TU�nvGTJ�p]1&AYbVQئp(��]�Ko�_�s`(�t�+=�pF�J����6^�k����eV_��k�]�jL-GI���	3U0����t�2���y����.l��)27��g𠢙R�������ҹ-�=`."r)s�N��7}�%y�2�wI)�*����gc�L�����tQH���[x��'g��4�?՛y3K��l����sp�0c # ҍ��_����~�d�	���y�����C](��w���jsڗ	^tbm�G\r����b)�A\`��\Y1��
�?v;`*��JyeF�@L}��
�!���Gz�xT�6���s��D���ۑʩ�01>$�������z��}&	�t����fR<V`c�mB�5t������x_�g���m����˕�8b���v_�yP-�ʪ�&�W�#u��%��H�K�I_����+c37��~*:)C���WXI1���;U��K�1e����(e�|���a�Bs���Ŗ(�d%��7G����C��LrՐ�����p��OO����.="��vnc}���RA�{ڍB��]��#�u������$SmE�ҏ���@_p°@�ab_[aߢ���P,͜��Iƪ"(�LB�֙�ϡ��\�*8����6�kz��M���2t�>��-��.n������<F�-6���
"�����e裩t~�Z��H����>b�X�0��Vk�A	�}o��N�Q���<�<�]��,��HvP���K��j�#_	l��r뷑�>ό�>�>�Ϥ������$�9� W0�$��q�
�y��p�ҩ3���1�h�@�WX��'N�h�p�$$
�C���D�b��X��;�^�m}cٮ��*���_��R���Ԉ��$T����0�t���o��]j�)l�V�Ou�iT#&��&��֍��ǲ�J��Q�mc�K�H���9M֛M?��/f(4���(�u�S�3 <����P4G<�c/s����#6t<	E�h��ӯ����8O����\���2��q�e�X<`@�k�V�ζ4; f�ڰ�z�x�l���Co��|������\�q�ƯJ |G;n�H���>�Ֆ
�R��`w��m�&�=�T�ln�h#�������K*��/��pmH'������2uS��/V[��F4�?M(@~�G(���}����_v6l�e` �� �)Q���K�bd�.	hW
�J��B��-,Q����g�Xu��Pޏ�����W��ڝ�`��wZ=����i�Ԡ{B`�*��56YH�~,�a��g�=�����?�v`#ᬆq���
e{B\�Z�7Ck�*�FP&,u�g��]� �xD8aƑ�5��h!��s!0�G��qFj"�س����:A��~�"�0��LXK��j3�Q�*�|!���O�ɘn�E�af"�}�}��<X2�͹����D_>��3i{'�H	���X$��AKr�&�k��L�>i�;��ų?��q86���"����X�=>kݬؼ��R)Q��N��$�d=8a7o̰����mdga>G���ϱBl�kd����"���E8����ufj�^�=��8��%k�^���^�	�j��X"����˥��	6���r�.��P.���i_����f�붣(K��x�U�`�$����Դ3j�'|c�1]�c�?��+��6b�҅M�i\�m�-_�>�}��(�HS�g�%4��'}�r&L��*�-�.
(noE爖 ?#��ë�R;�6[�d�o��TS!�q�N1����F"F"��v�j���8���J�tf���D��	��M��$9\g��JX3d�I\��ڲ�,pۿ�'jB�s���_�P3T���1e� ��h��"e���s��8�P�����#��Ѐp�4�A)}q����^��������D�e��F�nI�c|�쳉o*{�4�f�T�,�D��G%P1�I_���TXx��bí�BGQ-��[5�h���R�L�cR�
�$.���Cr_F���1��v���"o�r�S �_�� ��D�Ĩ���f�^� ���ۡNvo� H$!�L�hìVjѭ$�+�~L�
��	`�65|�_1��_�*�n�EM҆w�(!��o.��܎���~�������������|(���/����.x�)�|H�x9>�����R��q��!�+���W��v�h*�MM�h>�!c��.�N�"M��w�an��ۗ��{����d��S�����/:�(h�aW���R�C|�Y)���W��]�h£����RKQ����G�Ə���"�ݽ%FQ�C|{�mLQ�X��?�>��o�ăB�E0C}�+~���t��ܓrM(��m��=�CWdɸw�P��3!58Jԡ�(Bˤ�8����<n)��/RJ��_��[�������D�wLݨ�S�Z����z[ҢW��Nb�q���tb��RQ 4&.�S�I���t��N�'��Z775D#��d���;(���J{$�x&���;f�����J�KW��Ok�kfq^�|k�e��@�C���S(�%✾gŠ��$^rF��D����{�x�o^V�F���P����`qW|̐�$>����7؏0��S��F)�`k� `�_����A���Iw��Ĥ�h,�ŋv�xhh�B ���P��ְ��-)�>WA�޴�6�K��"很+�d���(��X=�T���v:S��%Z��7��8���^4sW�y/q��2�>=�?uW����@�5��2?>5�H�w��7&�G��3�c,��zM����#:�4�,eX{������$����5��4��U[b����+�i[6W��Udxy���.�Š���ȑ+%��z%"{ 
��^m�sJ`-5pr�%�`�q���X�8.�������j�uN��w���z���5�kc~'�����N�k�/m0�a�O7�
k��L^�coHQł#ж��0k&���
�G���w��)w5o�f�I�G%�Q/Ѩ�"jfF������z�x�N(�!^�]$X�(;�v
�5w�o�S:tG�2`������EB�@ߵn�����(�.���U��2t�-G�qj�q�Xq��'v&�p�����C1h�����O�/~4*�<(�ؾ�E�?絶"����ύ&�T�$�#;TqZ^���;���8�����:�v�f��L���a�/V��5�/��D���Wt/���@�1o�e؀1�n����"����l�O���&K#:9�YF��f=�����J>���i�f�˻��::���'�SS ��Hԏє��hB.V��^�f�y�����n_(�rY�Bs?#a����PT���4/"5#M���]0XG>İ� �R�H�M&$��ū
�FK���OB��Ji�t�p4�7h�ލ+1���`�6|ꉴ�BP2m��څ]m����]L���������K��n�w������£�jfm^AT�|S�J4hкv�ӐK�m(�����?���u��K��m'������RSh��R%8W����W���2��{g"�, ���a�wk��k�x74���a9`���R�H�,Y{�|���G ���`8iUԫ�VH0���M����O��� �WB��Ȟ.��zt��eo�>�M�b`r����W"zI]'�R�Y������w����2�B��Óڐ��W�{�\ivyWH;�R/sv|Zs�E���WHUe��A��O�J1�V�=��
�LG~$i��w�i����&�{��s��zԩ()h��C���J/�� ǰ��#hx�VG���>ǰX �X��&3b�:>���b��ϫ1Sjc�B+z� .�F��&���&tO��"���5�j��W,h��A�ܾ!��S�"ՑN��`����	i�F��s+��-����uS�P�ձu�=|lb߇�N�uF��Ձ6�T���A��g0ap[֭xw�?;���?Gr�]P�j�.�Or�R\-��!r�E)�b��M9�]=$
3���a�&��e����ɬ��+՚�h �T�>Dз��<c�I������*���Z�_^mt�:�v��5�d���t����,RJ�BH��;���2t�J�������7��d�gm&����m�K^/�8F�Z�H�c����B8`9�)]�z�Գ<Qé�:�r}��F����MTkj�[	Y�="X��}g��'�a������������w� �����-���æ���S�
���/�-J�i��@|b��Rd6F���a=^ɴ���1����$��zK�b����