��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&r�F���oh���ཌP��ЪV��2� Vvf�����jص^M�c��I��﷟i
�.�����H����P��c�b���&0!��}�N\�Q���<����f�2�H$���G��v��H���L;�՗���#�K	C� qH܉��e����'�ʾ�B��9�Z���l֕�F	��}��)�!<����j%]�%��i�WL���n=u�f����۠�\�?�Ǎp#d�C���Z�w�m2 HN��N��*=���X��|����W&��A����eI"��P�0�R�j�	+��JE^p&o���!V�x�����[p�%d���Ŕ�hv�ԈY�����%�ݿ��>��:8�kk�ô�c�
�ۼ��'��&����J[�(��g"`�fn�fTz�:t����)j��_��tv�t�я���L?M ¾�e}s���Ӵ � �.��z�Q�Z�\V�t?R��5�+��S�12	���F�77Y�1���C�A4�d�A�W�H�8�v���-��A5���L��ƨ��jl���3�܁L�����uV���?WO���:o�c W�. ���<Y�t�L�3���w� ��y��>�-�0��}Z��<X�*�͘��}B��o�;����?�Ѝ���R����c~	X���77F���<�3cMH����S��;��!W4ս�{��怬�����g��X�\&�/W��?�u�g����lR�7z	~'�����ѳ����N���D��塨f��T ����#�B�^���s��k�HK�-�Z�I1�4K�h	7�F��Ѥ����Xi��2���e�e����#E�� ���u?(���*�-beA8�]wk�a��A�i)��y�I;d����<(Ge����b��d}�B�)�/i=i(���4��0���Y�ٰ���a�8�z>d>��!�h��l��z�)q��pD�b#%#b��*|�t�B?�C�C�yE�]I�_]�f>��òa;Qՙy�s���)P_y���j�|�+e"Uu�V�[���ܙ�]���OQ��-��;��YOϿ�f)�����b$�RǾ06R1��O4�|t/�_�nսs�s>M�le������`�.EUMx� 6��Õ���-'���X9ArM�^#�c�\,GK`��r8F�fL%@��|U��0J�@L2"}ے�$��"mO	��L|�?�1O�9��w4��w�l��įڟ��H�$U�[m[�	v�:y�C�'��\�b�TR̮g{�:n`�z�5P�@ �"�V&�Ą����T�[��B�Ě�5��n��3�15�9oW����<�Zxy[�Ɯ����|�������1��/ �\���H���ܳ{ظްhH��(���eR~TGN4*؊m(��"��lu���z�VrZ��:��H��[H���շ��Z��Y[ˁtg;�/�Nn�U/�C��_x���;�v+���7�J�°�F�5�Z��ψ�nǐ�����pQ!?�6�M����.��c��Xx�Z �Ԥ1x�����6S�p��1�$ܧ�r���c<x��6��@;�@��}�@Ew�Il��_����-ީC�0�I�[�"�ϱB���SX�.�rlHieJ��@}(��B�kߛ
q[0�S�N�bݠ�ŇG�0��ڮ���!Xtk����D��:~�4���P-�s�}*53b�6h
��̙�Me���1p���Μ�Ӵ.8���:h0mK�f2p��E�?�@�q&
�O�����sD�����ʢ�T�-�X��X�"!��#37/�j�c�F8��ꡪ$�� ���-�����x��ܯ!�^9����}Wq3'��IK�.Z���//��6)t����
Y/xבșJ1�&��*��aR$@������,�S�� �B�-e�^j')E�&(F[����Yd<��'_���U�J���_�q��T
'Ɨ�^*|.grԵ��a�6�i�˖^CA�>�+�>f��Eo-3 2V�D�{ܿ�bᄑ�K^^�&,|6w��H����x{x��[p��G�ҏs���_n� q� ~��X�ߗ�e��՚w'�I)Yo­��?z�:@�|(�����`��vs���.�PP ���������ov�y`v�x�΍
|	v��U�
d"��)J�2͑���i�_"��^�IjL`ڒ�W6V3�P���!I �v���