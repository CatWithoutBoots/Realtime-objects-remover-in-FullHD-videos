��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&��^L�h�m��uXҰ<.`D�iL[u%y��{����|��G��u�e~fc�b����K�z##u�9)�_+x�s�{������p��8�c���7�"�4H#���;������l�k�p *��o�G�G�&�]
�_ƅr��ЉJ�6��|.�Z-�}!�#�ձfE����H��=]#�MB[V��J$��'��X ��RS�Q���1M�ն��$���L W�����@Y�֭�
w�39h�J6���xI�`�US�0�M���$UX��(�P��������������P�`ⱓ][����;b�Bw�6J�&��"m�6�>eR}l��q�d`�e<��3z�x(�z��)i,q΅�t!�t��:z�L(��ח\�k��M ��A��=�!
���/�_G���3��<3�����u���T�lϰ8�-�ؓ��<�g�L�ȪقG/��
'��am�+S�%B��������7&��*Q}S��\R;I_(��/�n�cC��q��#���N53�^����
`���f^�Z"�-�޳��bwϖ�
r���N������T�����D����h`w^gV�-0���4�v5�a�OH������Q
[�}ȫ��j t��,�B���qD>��&�T/�^J(�Di����z�E	En�@�1�ːdl�m��5���՗�g��ov��a���*�!����ZZX�d¥f�g}=��-�q%l�A��8�\6 hi"�_�Y������y�f���]��BAK�랕-�=�h�\�5ªoeZ6f+���L}� ��F��y$h8��ӱ��f.J��s��oǖ�ɡ��{�yQ�U�!x_��9�'[/����.��~*dA�����Gr��췝yaty��9����0� ��ά^էh+�ŕ	�ͻl�/ ���|��+��0�JP91;���zc�v�(^l&BDr|����Q\IE��2CΌ<���� �#@���*��b��������
����~�>ԣݔ�=�g�� ��-��X�,�`3�1
7�n�mp���Ʀ1O�1�Ze/����h�S/���ͅ�57���,([΁��6�m�*^\Խ��o��<�~"e�]�6n3�"�%YrHI��*5��S�C��0z�m�/���vlJ�n�F䷯dWҶ՗�����Vt��������t���
-AW^�j�Oz�f��i{S�g:}��1������9!��ݤkU��-����υW�$n��.�P��D���3�g���#}�C~)�r�]�hln'g��܅Ϳ���N��� /׌��{놽��@���7˘C�&0��o�gg���	��A
]3�QCm�"�"qa�/>w<A88c ʬ��?T�MJ�4�ջ+le��4��=.�$'NRU阀�*��l��'���YS͊ů��<�"[!�'��˄�xQ��4�fU���'�e>�TÙ���ռʥvX�wTҾ��`��*��Y���S���uI�-aG��N�[Iϰ���<.�M>,�|pz���\Šd?t���zH�<�%,�u�b�j�T��_�i��H��X��Wi����vz�Ӱ�l�n����&9XS~�Ų�q<���̒�h���i�jg�T-�����݌��牘�A�����?�5�x�}�8S��cn,o�&FU�u�e4��Lm�si�k�����po#�A]�~G_�L7���]7@*aR�OnVv�][�]
���r��B�
�'�L��������D׎�pؙ��]M1z�"���{@��V�?������ hRz�o�J�:}��"I�2gW�8�
w���'�B?��Ѯ������m�6��6�[_tкr��QK�|I�/��x�|�嵤u�����G�ǁ3I����N��j�j�IB{E���ӥ�2	 �}9��0�*�>��>fk���iw��TKU�5��@�q�*E�Q���a��>�n�y�ew�l�v�B�=�e�\Ax��;,�*t���|,�<-��m�M�/��������R�p����ѷ�UԼ<l�A��u�ѽ jF�Rj��Q�qZ)�S��&�\�[T�d��`sW"�ZuGg��׹( !�`���!Z�B ��\��ͅ	�`��m��(��t�(o �=�!
��_�Yw[��K���n���mڗ�`���!T5�˚�8�VT��7�c�U���P�2�]"�$�*[�y�O�Oi1�x��ki�x�n����R��/�\@�=7���R~����=�B����B�����)U#�W�(��/d��(���g��$�%������`B�A��u����NuZ;�154�I(�q�@Д�����Ƈ�AM/�ԏ�@���l
Ja��lg�3j�c����O��{�=�DV��O6���ȥ�i�Y�XJ��f=�;-� �k��{�ᕏ���߮��N1O��ʎ���+��q�O�>�&�8��^��J�RgLp׷5��I�D:3:-Qɭ�uo,!�2�xk#�D�(�;ф�� �O#��|H�ȿ�;�Sg4q�����pR@dN(�`�K��O9��X'7ɲ�u�1B�i�gr�]ӅQA�foF��3U~��5xJu8�1���}Q%�y�pq�o+IJ����`�=>@xFa�^��af��l��3@#8���W#�_��)��������m����� �q��Ό4%�a��ւ�:���:�� �Cg(�!�#�ת���\&�[��֮��%eg�9�Vo�C3�$uC��=��˨r���S%�W+��҅T��W��E� �z.X�B7�M@}�����.s ������~�ٱ�(��V! ��R�Fz|%�6^M��E�u,��8ѓ#X������mG��ܘ�\Ջ��!?����чb��vm�8y� ���J9��Fz?̢�U����^�~V�9oG�#�K8G<j�Q�Dr2�6K�a���ISh\�S2��'�qS�>�]z���g��@���,��(� ���)>��a.)-�K(����4�&{�\�$�g�;y�`^tӌ����U}�����@g9!6Љi�I��Ԫvҝ%6��k6����T{V���E���Sf��;snGB2�Q������ 7�����}G0��WqU"�tv���UF@Etp�
���\�M�<�4��_z.J���cDm�U���c� �LR�jO��<e�wj��PM�� n7����kR�M��S��}PL��9����3����H<b�;xǈJG6��#�~�J�ht�}�q-�ʮԥӺ:uH	0���/���ob!�A�J��0C��}�I�i�R>$t��r̽B�/ �4?`tI6�I�2CK����w�C�n�� �ϝ"��ϖ�'���\^��4^�|L�HCVAd����.�U�F��V^8dX�)�'m�34E9��5Q�&Ļj�%�W]�m�x}i��w��o5��L~/pQE�I0�ΙDg	��V��2�s	ۗ�]��dE�JO�]tW8v"���W䱥*!�u샤{u���j��|S�M�Ѓ4�k��@l�v��$����_����N6�E?��6P,��Z�9t�W�i!u)���꒒k�0+QS�4�4 �%���l\N,�X-N��$i"fq�T㟱�1�i����yx�	!Wҕ��7�v��C0�2v����[=��N��9�a���fzU�	�bBf24��¿��xY]� �k1�`v�3<F3��J?F�.�����>����_B�����+�

	��� c~n�P�@��ߟ�]-�	�zu�[I�QY�h6Q�X%�E8j	�9�:R�^E�/�����E�	ȅ��0N���fL�Wǉ>�N<��R��L�P`�GM�٥M^�d��A4��ر��Y�i��*{y-����0�%����jK/Ye������d�k��Ʉi��>��_�������lI<M���<î0UЙ]��)7ȓ�琍O��ǀ����(j թ�_�*��L�kJ5�K�^�74�����1n�[��`������q�R�
껠!�������84�Py'i�P3�6^��D�~uɒJ;85 HSL��ў�I��Z ���յ�i?�(�O{��ޯy��g����A�n�kJL=h��6C��0:�6�K�g���Ǽ��Oh�����9`��J�Dlh�)%%�_e��8"�I�?jU�=�|�f�e���޽�o���a����@��;�a�,ܜ�[�e�;9��Mh�3[�(�>��&&�J�����ɝ�.뒶��m9cx)�l�~�S��x�0L�+yk����A?h��#ȃ�5��ڏK(߭�C�|dr/�dt ve�I3��1�^�U��m�0�)��voV����b�DL�l��Y�;0��P<y�Ȑ<��O^�.1LS�ې��1v�� ���Z}��K6�K�hB�Q�4���Z��X�bS�z�m^�`�"ј{�P>�.�t��
1�|���R\��9��t���Hi����Vt��s2�l���|��$Od�Q�q-��ܱ�n6���5S\)��_����*���i���OLO,����.�����Ddo+�鉷8�RX\�]�e/Z�Y�!�\�gu�AD��N
Cޱ�����Y�)�<�	b]Vۆ�R9��.�.�-ϻx���P{B�]�MaL���#ytU�֤$�UZMR�~#������#���෮��a\�0���Ill�������ߚ��뀃&#t�?7?0@��X��K��h���X+���cz��q<A�m
B~��Fۉ�O\�ť��R� x�h���~�2h��)7�c�?����nga�1��|��Y�d�v4lf��;ό4�ش$0|w�Iu
�_�����{i�(0<?tv��z�@/�>��z����	2�Xd�?�%�m�1��7�ͷ�b���W?���ҏ�/[��y�%u
��QY�I��9n����9��6u~�R��E	b�d��? ��H��(��0tI�.B$KC�t����\���l~^�$T�˓G/c8������/�|Y��{&1�������C�e�
~��/֠��@��p�G��͒F�=�)�U��'�qƊ�+^�`� �bj���`wcϤ��>������`"~�&Xf�Sqfھ�gQŀ���'�@�V���S��a�w9���ރ�O�o��j�E�S3�v�P�Q�
\B;?�q>��c]�LN��;��zJ7��{��x"t��@
�)
"�_u�����ٌ����:�W�dn��L|���{p�8B'��n�U3j����vu�Dԝӄ�~��O��>0�>L_7޿Țoj�,Ѫ����Y��s/?�e����Oqu��x�;���"�0,�4�����F���^y��3�e]�AJ��!WBd�F�a�!�Ǖ�%uҦ{�<˂����P����&���#֙Ӌ+s����A��dw ������J2<���zwS(F��೭ ��P����/r����9q6���^����F4��ut"���X�f�����5Ay���$\��E�>�]Z�BW#��I��iu2�c����� �α
c�mț��`�^�ț�D��������������݇.v�΀8��\ò�YRl�̸��z�%�dp�O������=��2�VL��� l�M�/\�2yE��1nʿp�
xtë<�����I[2�r+��2B1����m��j�<����S3�ጫL�R��9�#c,����nM�3jI$X-Z�mã����C��/�P��G[��qf���>�Ŋ��[��j[)����ya��M�Re���O;�X��넯�DPBU��|`�I9�,�gD~1l?S��_��a�ְ�\���a�"��Hn�r������3Joy�1}��J��U��%���$�iP�����QӠ��R�7Gh�Zx�0�;<�҈<k4Uh�p*  r}<8�z�1��[�Ҹ�,�߶ +�:{X$]�AQ�!X�zui�+�훘"���ȩ�S͚4Fl)L��竟c�:�=��=X���t��a�v:����f�j���@Q���/�p��� �dZ`I~�x�Uxa��"�'w�rp�FA����:i���	B3������nm����	��}_�Q��4ͧ�9+��-�dBqC\k
�.ȗ�1H����F6_���*d�'��S����`��_�t]�Y\
Y�/���Ly���3l}�d�����o�c�\�>#=���]�-ۄ '>s��[������) Þ����f
�y�\��#�[�&���ʸm��'T�B ��V��S�� H1��4!�@��Ԁ���YW~vɕ�d���n����7� >4��F�T���o�����Tf钣�y��OS���p��|6'c7���d屴�xP��y�[��\�c��T@i<q��l�J-��k�q2�n�G���젲	�׮W$�rE��N�R���*~t�������%�\^~�*R�I�j��u��hC�}��u����YY�ޠa$��n���Ē�N,)�T@��.n�뙽V�x?ݝ�<�4vW鸈�R�mo
�h�����` �h'm�ȣ�v�up�̘�&�xx1fijB�+�e�yk�CPxh�[إ�pk 	Ѭ�i�)�H = 5�����58�[_�n�;d'o����pzu���,1������Jo��v�F߼�u�޸Bp{T) �\r{�mq�*��V#Ij}	�(R��7��-v�Z���~�Ϯ��?��0k�ڲ|`z�9������~ߚ�i�<D@!�U4JP-��ĪX���Ӏf�q��Ҧ�������4WlS:;KZ�̸F�/\�b4탢�z�����6�wB|��!�Q��3�j�F�G����v�x�~�;\5�F`bȔ�I.:��h������N1%���{�8�gLK?��z�+��� Y�%=E[��[��p���� dkrQ-@x�*�o�BN�����,e�D[��H����i�-�,cU����Xć�� #�0�vx}gN�e;,���(�����
��ӌ��'u����>�V�q���a�k��4���;��]��T�WӺ>��B(�5�>y�,x��E��7U�"PW���x�@����BGh�EE�s-�6XEA��ԠRkQ0@Bm46�`	�Q0��i[�<_�;/�[�]���D_ ��3UH�|p���4�nZ"��i������r˗k�۱���$m���@{�M$_��T�o��H�}���^~�C�"�8����E��gz�ɱ[��wH� �)��m��QA|��o�h��@~d��b��s��"-P>����e� o�,ʇѸ{�A�s�*$ $9�;T�$B�x�_��CK��g�![$�h���Eܿ�<"���|���%�V_�w$q
uz[~�\ �m!fS�K���8eB�~�9��E ukS:�f�2��
�������r#��N����t
�������w���Ya����BhC�e���W�eP#iOO3�\bϸ�m�/�xA;�"J�<��A����-���}��XHK|��x������[�Ƿ�N�!�s���������t2{c̡)�Q_��˝%z�1eX߱��!թ�k�r�H��cF���_itk= Q��\]Di���>�r�z�?$�U�����Sܫ]��iu�?���V��H�`&�cӸ,� �$��C.@ϓ���b9��b�V6�i.&9iB'����t��mJ���"��o����<4@��;}��W��Ԡ���?�I�[@dCOP�ɝ������s�>�S�b�vK]�@�65nbJ~�4 3�)����]%�y@qC�J�����&N��se�x$��q��z�f�����'�l��p4�3�V�fG�.lPrѴѠ�]GĹ�s,%ZB _�$2��]
�bH�uxś�P�>޲� P���p�������+D0�~e�*�j��8���;��T�$~��N�-��*�Lb`�]5ݢ#����*�@��i�n�I4�/C��d�W�&,�qw��$1Z;]���6�CEu�M��zY��`)�+�������0O�W~(�_z:���!��Z*|�%��6�ڀ��˰������߲˵�m�w�ni�/>l��ҧeNx�+{�Y��%A�΍M��!��<�Q�z����x���7K����c��rG�sI9ߌH����ϭ�3ˌX�蚴�K\O��y8�R8�H*�U�j<;5[`���\�-N��<�U]�l_���1��Z���U�*�?lz��@�N3��j� �^8� ��Q9���ޖn�3�1SeQ��χ��M�Ѽ�O���6�Ժ$�}���:3I�
+���*5<,dwO�`4�w���nhݮ�A��y���vښ^����+ۃ#3E�͔9sǗ�/�6g�@�n�����FȆ8qF�t�;�І�:o��[�O_A�����:Pbev�.�����t�A��q�Q��ݾ��F���{���� 1:�: ��2��k5�$�����\OH(1���	ִ�ps��AJv)n��f+�]/g~qp����5/�-�Xa���	oU{���H��˃���l����I�_ R�PT�+�~g�(��S���XA�'�����P{����?O���ڕ0N':�`MVǷɀ{ЗhEؿy�a�y�\/�E��Ƅq6�7ƕZ���֍0ǵ3���l`}͕�����i������Ms�GM�@*у�I,��ӂ.g��$���;�L?�(�������7Q���4Ŝ쌻-��l�I/ν��qA�v���aB��[�`�ƈ�Yd*��@ pg�������3�X���wLܕ5�?���8����ҕFDt�w�mh��2���Thޚ��^6$�t��z%c������%�xږ^�n��/�k�:V�ϳTv��Vv�4Um
��*yg�Ս� ��<�sT`��2o��Kd�<�r+!���к�ʥ,�Z��P)734��*u�_�sy�1�_m\����_V�X	:��ğ����r�+�/��bYeU�c{WLM�zoG{7f�F�Z\!i�����@���9X��G��ubV�n$_����D��)���=�Ø�IhwR��C�G�0����S��-�	 3��x���Z�	3w:�:;|H$@��-�Y;�Wb�ɏ����o1�w�h�vN���|@-��E�(
��ؼ�]�(Ǘ��z�a���g@8y����=�v,�ON`v $/_��������m���	6�)t��r���x~��yZ�n=�Ό��Gܿ ���u��ҷ��`Ŷ�����g�ȧx��Qӽ3lƦ;\�����[
Z"후�+ݠ:L�?N������Do.cR�\�:����F'�;H�{}��%�Qx��J�[C�!&�P���=)JJ?�[ˊ�ܗ�~����ُ,JA�$�u�(�%� =��I�d\`4G��J�p��\�T�b����Zr��80`Q�ח�?r�4iI�ӑ {�9he0h�i�6tU&kQ�	mK��)4��e)��J�Ղ05|^��۫3j��$�i����!k�mVi�B)��9�#$@4J&k�@��p)�h\@����-�auJGspD!�����'�: U�	���	\Ϸ
ԗ��h�H�{��O���ߦEf�)5�Ua�9@�SN	Z)��ſ�i��j�aޘlP�D�x��K�iҾ�#�lXP���.���Y�ZJ����V�ps!��Ed�n�?�;(����V餚�o&z�����r�R$x',ǚ�<dP56��p�p�&��}�r'W��H8�z������XJ$!�d����T9Z��)���_ ��ǅ�	&Չ+*��;�yS2.	]\1�h�U 1ՌK�]+�3T�@��Q��+�C*݉��R���M�>+������:,���(@!��2ɹ�ԅLi,�e���L�H��aL�{J����O�8�Œ�E�E�pX�c��ЧFG|��Cֹ�y�0,�22�W�흵U�C@�w���P%��<�$fO��<�����|V�y�rO���\�^��F���x�؆�N��#������H��?G�^���9`=��-��l�:���b����"��Vc��$���ukWa��(���,��R��;������i(�U���S_��f\���/��ރ�l��ҕ$��	!�(2�����Hl�o��}̅Sx(j��-OЏ�4�}e�9f&/���oc\��I�R�<m��P��3�˸�D��ѾQ���R6%�(�J�'�,�D��Zu_����R���ω=��	�Ί;���d=��Fa��� �;#\��	��M�x�$Jo�f�A\_pM�*u|j4}��S�ͷ��z�̆�c=o��kG���΅8�\�A���5&�=�k�)MȦ�ʻ���z\��r ���dJD�T��LF,h�uO��ĝU)��WN���a�{7�ڃ�e��!3I���,���;++�j?07>"��0��cPLKT���+T��@Ķ[����@\c����X����JF�w~~N���<l����<�}+�V�_r;%��ތE�,W��йg[&��6������#%��ķ�-2O�X!�]��y��I�5�����>Onh$2��0�T!M�ӖUɏd��va�'�<#����}�|�X)A�]���J��	�0����A�
��X;�~ ��UcŢȖ����"��n�D����&T�s}���x�=J���欙j��Y��2|H�0P[��5����M]=Dn�D 	�§)�!�ύh�� ��&1?�k�4����".bv"��F	<�}&p��>DY�a �����.�I��f����Y!_���ͯ�vŽ��������j`�*�L��˃+�v���kL0j ݧ��l�>�gF���~��^���xx8Uj���=�����φXN8T����RNnr�=���L��W��)��"������/�����K��C��W�Sn�ݘ�}�VC-����B���7uI�����5$5���փ_�c,?�^�m�Eʮ��v𴣰�a��D>��Jk?�,gmU�C�rd�l2��J��P��$��9	��"��b%��@�ꢼ�_��~n2�I�H�,'=LP�Ks�J>#�e2�'�#e�t�۠��x���[�T�5����OS�������g.aD|����:��HQ�0+Gw|�&�l�I)5�b8��dAC4�G{�ܓd�������T���\2����I��D4PQ����p��yA���_g�z�1�V����-��%�)J�鑉�"���=��`-:�Vk�T�u�"!~j���YH�p��[/��LK����q�@�Nc��$�(�,�Z���[���Ąi�G�>v/�v{�丌^�m $�M���A+�>	v�%[�L~ɾ�/f[K��������<�~u�QF���_/A�����5��ns�Z�;.#J�O�P��P-+f�z:���co�9��PuF�U�ú?
c�Cm�&��,1�T2b�P
ꐚ)�Qp���W�O�N��/g�ֺ�9-ҿ��[���EK�oS�bXT>��XJ�k�T��ݼn�U�P��N�f��<��_3�����ц���/���c5��zsٕD���VAJű�r< �,Z�HA�@U���#$OZՀ�	��E�<b�=�#�(^�l��Dc��X�96�qx�# 'qC/�^���)p�-���{b����p	�#�/C@�i��(�3��oDo�Z� )b�<���+���Q(:R偙�uUF���9�Wt�C�w[tJoP;t�Zp���Z��fO 6�6E�82o�[��]�����XkB��b�'��Q"Q������o�x��7�� �a6�j��w�6�<�bJ���XTN�0!�����u�w��Q/����<hKMўcW;��1�v0�?<��#2���w��c�7h�L�M�`�41�M�����ၒ���.aޫ�.[Ͳ�� ��֤+~��|�#/ �K��!.�A׎ʌ%��G������ ��"N&'@��y=X��>h�&3E\������	Z��ȏN ���F<\;�K��/�8���+Bd��b�)��y������R�e�)NJ�_�V��[�W/��+�)����um��}6�F4>��Y�K�ȥnuX�O�o�L�}���u���Aǽ��iؖ�3���&FP�?�fGw.jw�:u�;����&?'�~>�A���x��I�Uw	�o���񐭚�U��W��?W`��3xh.���B\���w�n����A�I�����1z; ��� �_5��|w:�}�n�P��{/�Z�Ֆ���|��X��Ќ��e?dፃD(��4uBj4QU;6r�ݪ�7�w1q%�z��Z�A'��,��ҳ�~-ew��E+��*���HS�=�/o��K/l�,\�|��[�x��G�h�����!;�sV��y�I�,��8�r�Z�"���M*�h���#�tv5�ҹ@���0oe�/S��Y�@U�-`}�'�-UЮ�y�bf[d���t����W>��i�~Ng4�g�g�c�_zM֫}�'�����%Jyq��~��M��hT�h R. �<s͖W�AЬ��U�����5x�岁�+�� ^�L%@�� ℓ4ƌ�t�����iJ�AH�@}�"й��疕�{ʬͮ���э�آ�\l�QΘ:0������c��'���>��}�8ג�R-U
 5�ޢ��h��:�gx�-Ĭ�3�%�]��SÐ�^}Pr��
k�%c��'l�|�Y;��(�����̿y�5���<#a�)!����9ꍪ�:aU��f�¶z�P�?�i�|�#װ
�T�|��4��r�~uZ`&���@k�,Ч6f0ʴE��������&/g=���n�]:�]�cH^H���Ł;�!�{���~ͷ����1��yK�$���0��h�H�<���K���"gO�I����􎢬����={^�KfX8*y�$e�:T��**�f�q�a'�UKｰ5�Hi܃�\�;F���VB���ꍔ�j��G��ʰ,\,J���P�n��I�1�h�va^4�9��\"}N��M��Zlf
/ߞ�\��u�T�y�	��P�[m7�=8��|�z�i<��������o��-���_�JJ:ɽ�/���Z���܍{��{Z�̷W$ ��/����j#Ư��k��?�<ƻ�ha�U�9�7|��n[��Ȍ0���԰�7�&5�@>F�ح�5U&���(���U)Q�϶�=1	wm���5��*r!2K��@ve9*�v�����@d��I���_@[������`��3H'ҝ�&-�y5m&𵑙�j.(.>	ĽPSʅ(OeR7\�܄������<�j$>�l ����Y��hoܽZ�go�[����5���W`l�W���Yd4���j�B`��� 7ɠ�n���%����9�0�#-M厨REG�i�g/�v�p�U;��Y3q���.��5���#�U��,�����`����\yXo�D���Q���X��8%���E0%qAW���� �`���4�DK3���XI[�j�s�x0��p��-�2��9���G��yqk�b��oUl��wL#�D��*�	��{#x$�y�� �*ll���P�m}Y$R��z�k�8��`Chsr�����y$Lߺ�	��>����T��j���5�����g4{ld�y8���� `'R���<��{O����Ge�W1o-��gLV�(�1��0�� W?�7���>j8C�0��J���f��B��t5La��;�l�܌���Z���v�͎a�Z��<߹52U'����K���4o�
��O�X!&5n�ƫ(D�;���S%�Aن6KI�o��Ѽ��
`>@~?�]���MT ���F�"�ط����^ yJ����eq��a����E ����m�"������|s����gT8>�tݭI�]1�dl#��;~����;W�x��gph�k.��V�K���m�y?s�\Gļ"��Ll�%��bv�}�χ����E�5�1]�w�Ԅ���O\�%a�.�݆�����M����޺W���3�
auW���n�I��V��F����Nt���2DoId�����Q�5h>�_��ޝ��eF���1��i��� ͘0��x��$.U�c_c�r�f"�'	������L��#&���T�
�>���Ǜ0�Ϲ�D̇0q�tk��P�P8`�(����|��@~���e�팇��1��aR��P�\�D�q}���D���0	����j��Yk�U/�f�'�4��X�|CmXOV��78&�����)�C���',8��W`���6on�)b2�R'��LQ�ԲK�=�����Tfb�>��Eb8],5xA��
��`�'�G�yt2ؗ=��f�o�_Q]�Nj�WQJ����h�n)�A��� ����}�RH��7s�M��RZ�"G�ӈr�\�5@sx�sQ9R�sR����<UNm�za����W#�og&=�Q��K��8a�:�e�X�N3g�w���M~%����LFM�J\9H��3��x	��#�<ʛN	BA��g(���7A����ɉ۔����$��j�(��Nd�q�}��]��������3�xS��#5C�D�"]xvH��4�,x��XVl~c>L:�Um��Ad������E����<MJ�%ƅ�̹*�*L��� l�m@.�2�b���p�Mm�7M��u�U�e&��0������y�M͙U����#+�J^�Q�PUs�q*�ۓ�3�drH�����ɡǣo(Og�.J�/��ou�;�Q���,l�_�f .�ޜp��m��nEL�sī<$�|�m�~���Z�P��
9t�y�&U��}l���H���HW�Ï��>�8��n��UY>>-��R?��zU[_�I΋��]��Ǚ�/�p�A�;Vk� �D_�g���q��*��M�,�]���<K�7>E���J��QY�8�w�0h�ߜ��t8��CZ1��l�S���9�5�k��R��Nm-#�up�Ͻ�tx�g�{'�R,���������Ek���
y��#�E玢�}� $^U��$�r(KɅA��\@�"A��+�|�j���e~c��VM8#E	Olj:H�&�o�}�F�S&�Ul���T4�NL�C� �	�ȢN"H%Cԝ��Qz1�7��q���ۅs��j�da�e�� k@�P��a����5)Q0�-RPs&�������[/.6�`�3�{c��n�/r��X��B�[p�OB�oXh/����,"Cm��Á�+*T�;
����+"g��~��cҳ����,0�pl�!Vi,w�f��	�nt~(�b�x]��xI���t^���E�Q���Q�R�:��O�Q��塚�pũ��!Ij�;� #RV�Z�
;�l&�)|4|�	r�Fd1��|���d����9BH�ltçB�C�b���OD*1J��M�j�7 Klx]E����
���KG�N}f��K��1�A롽��M	�������߂�\���@�-�(o�©.�j��-��Sk�4x���������/}e8�VB���[�}J]^T����a_�ȩűTyk�Z�m�M�+m�M8�o�{�#i�]������^�V��6�״?�k���'4���c4��Ϫ��ؾ�����F>%����S�d/c�H��C������6��F�M��I�P'��@+3;���c}X!��Ю��Oץg��I�k���:�j��0��4�r�k62$���	cV������>/��"N�Q �p�ӒL���nQY?���̮�����v�9�n�OS��n#��)�Kjjϻ�s�PkE��]RmؚvQu?�����F�G4L�m_佇�(:��.o��+���@�h�M�]bS.�u8}�����D�$��&��T��XŐG���[C��E.eyvB96d��#@����j��3r̢�*Y�`p�ˣ��7�Cc�Ys�oW��1��~-����V�+��ξ�d�yl\�!��?u�V[ke�!�_�ӏ��Z2��ϸ��o�l��u+�sm(֪ۮ�^`��Q|�oBI���JS����P?�L�V!f%o�P	���[Y�L��g�i?w\��$��{@(q�g�7��wʗ<�*�p|�%��D	�+���
�/c ���uv���M��w���T���\���wP���(��J¸Z&���[#X��N3m;{f-�S�K�����x���.osp�4��2�F}���-�,#��3�*D�����fl�*��r�2� ;D.�~�W��\�[�  �<r�b��ҕV#�ȺpTY��vp�93�_��Lc��~n�J����2�Y;6��ȵ,˚`���AT2�+->�PC�<�F�S��5�~�.�t2�k�e*���A����u3ٶFf�@���+sg�|��{��N**�E�jy��O�B=��oC�a��F�|��D@$�8���5U%�+-\�hv�L���E�ms�KmiP���4~�s[��&y(�M��O�&�{�vb�?8Bn����1
 �]5CrC�J�6�@�o��mz��բ��\�4��Q��x)L��uki�`��_0�N��ԍin/�'��::of�l�j�r�:��Lgã]yq|�����l�9Z�5�e�}t\���Z���UA���ݷ�����h%ﯫ��jT�*_�����l	.<�r��0��������܀ᶭ�J�[�*˙B:�ps��+����Ʃ�[oJY�����.�W@Kpb�����M��3U� ��:��8�Shf����j�ԍ��ޗ-��e��Y��F=!3p�>�0O�	}x^�=7P��BK<��@;>JwP�����">s���F��(� GY/l�!����bR����u��kBy�+Q4	?��D�Da{�͚4�<.J���z�E�7�.�moB�y�YN��E�5���S{�M~=��)��"Qc+"��Ը弓�K�zk�*��dY�M4�����y�aaI�)���iø�\<�Y(?�e�I��꙼��O������=�|iyI��C�>hDy(9��b�����hNWˤ����$s��c����*�+�)�I&�^�o S���
"1~Zv����𥉉e���R��,��o��ݺ����Dˋ�P����~�ˬ-� ���V�Kp㠔�粮֧�ӡ��h6F�X��T��z��&���.���dƂ��c���4�MZ.Ww\�X6�&Iuz�cz�0�~�(��5�\���"Xc=:�y�VbL�9�t��q���; қ%���π��"����2g63�,[��_OB����ENp���c���?���I
����i#�C��B:��7r18�ze!Ƥ{j`���`�]�����m���\k5˩�	��iƟ��E�g�7�$��i%(9�P���v�p@V2f�U��&5��`��VZoK��R�1N&+���)�b�Jw��d���O߽Cڠ��4�{�����B͊HA�Q�	JB�3��y�ɠ���>�T�7�3�9�4R��Fb��O��E�2�h�����X����Q���4��⎦v �B$�<ua8Uy7���a��}-��4oj�&���<I�&��#�����M�ʜ՝Iu���o�+�h��B��R5�����S� ���ɂ9�2�1��q���������.�Ȳ5*Y��5M߽������.:3�vUV�1�&l4f�܏&�_�[��aԂ#�ApǠ)����-�p�}�g+a; l����t�Ѵ���:��Uۊ�=I�|f߭�����z
Y�.�����˪�v��%ɱ���w>)\�nA�_]��Zd$Y�i�#��/����nV�RB,OA���P�\6^��/ViI�>*,뉔�ls���1��\n�s�,r"�i���l�2"lǌ,�ՠ�KoUǏ>��ß�Es��r��!���H�r�jwh`Gz?2h�`�!�a��N�dY-��_�׀D;Ƒ��6�� V�0g��M O�4�f�ȪF���|UÇ�c�q�B�3����pٯO��p��nOe��a�n#��3��-�y<s�wW̴�.�Y�Y�\���{��!�ᏁKr�w���������^+�:�<���(g�C���{xf򵗑� ������``��)��Y- h5>bSn("իZ��i
�5iQ�o�l�h$"��L�>'
b��C�44>�TZYE�O��4l��1s�9���|NN���c�(ێÈ�[�d~�+�o�����eI��,���yl����$�Bj>����5aY��\���N�R��	!�+	A
�gp�W������%�M�L`'��H���[�x~�S�E��+(#���v��|7P����.�ا(�	�c�U�Kaf�;Y�)����'W�����N"�r-�/M�0LG�L)�����x{L�g,R�84$��QL[��0y�������6���0 �y��|�W��,n� 6�z(��ڰ�w���4�+���w�y��1�۲k�Ͷ����#Jj)a���tJ��h�`&�!7o��Y����"��!�6q�YvS��`1�N �T�pm�Ĩr*6M��$���=�ٰq�|�u���,%I�i�v�?^���PE-�F���� )�E��$�������˵���
9���G��n|����D�+��M鵘w��Ey�������}����\{D\�����'a{
*���1Jlt�WF��a��ty��}3���xE�a�*����Uo���;�%e�A���̣�ENt����W��{��s�������p��jA�5M���[�r�i��X����k1�|�5AV�`2m�z��I?��P�N��U.��t����G�p���y�g��G����l1�&P�n�z� �Y�F�E�=�7�K�\	G��t��g�6{5ٔ���~@@��#�+�.�z���#��$i6)����ق�6��j��{�-Fޣ���9�����-T��rs��Jɭ�[�`�CL�N. �+L��2�I��=⦚��������nK��v���y�^_i;����p�٧�,A��TF�-�(��?��s6�N e�07,�^��ZQ/��"��Ïi�����p������7C:Gr�er����&ſ�u�1'�U�tei7��"=��m�p*0 h6F8D&�|�vu�BeV�y���P�aB;�_�~������]�]�����~5���J<
J��Ie�;L����!��o�i���G���>��"B���ZуktʹN���x�u���oP֦�܌a�'��$f��)�����	�\z�6s��kY�����/X��u)�0����.���m�U�z+���7�4�.ϵ�[���-�[��-�n�$֚�"�=�[�C���֏2��� ��'D��[Y3oi��4dڂx��"�����F����N}�#:�;{}!F9�K�U	����[HY�}�*X�'af����sE��g��PO�e��N������w�>tz�x�4=f��>t��K��e��9�ڥ�w����D����%��Zi�._�M�:�d���`JA�#Z�'S�,����_u�XD��kh,��>:.rE�L��d�4�l���,�ܞ�U[�7�%����`�.gr��'����i��0�"}C�t6m�A�N���Y�6v�Qʣ�3h<��w���*�:��W��J���N�� �������_}�Hx�����bHN[v�l[�:�����3�N�GdGuP8�����sf.��qFW���S�Zso�7\ը��_��� �}ޙ�e��4��8��c��WN)Whyv���[D;v�����*[��Ȏ��ĩ&^�[�B��+��(��/�ͥd�Ț2�Tq���j��br�w�G�C�=�f�3H"�ÉD./��Ȟ��|�N���h%.�PN[��c�|��s{4M%�����T4ґ�#�bL3jG@T����m�º9�%|FY	���lCͬ�:#'�p˚(�6|���Wv��g��˫�y�	��`=�"���O�%-��۩A��o��W�B$d�:�S��V�|���]c�	�_�Lt�˽���z�j�P��� ��Ĝ�l= ,7<T!R^�a!t�S��PU��)�ȿ�R�"��o�|R�.K�E�`I��LL��S�������=z��`����P�����@�X�@-�h��,[��\��';�$D���k�D:t�j�b�!%�W1��ݺ'�I����u�-b�B��{��2D>�^O��8����>�cW,W�����X܅7��@�hR����}Q�2�YM�2����\/�C��]��s���q,���_����H����FN�Z�R-�{����L������a�����ϛU��*�F_z������c���mгn�a����'�b���4��+ڥG%m����x�T�,*�a0��}�Ib���Fj�cG�6���D���"Ъ��+��H��Q�R��Ũ�y�5��g�"o*H��{~��ny� 
�`�c��/�_O��9,+��Ņu39�q˯[�dNH�U���Y�X��
vA��R�.e]����l��z�3�.����(��S��*��=U�q��-��N9��ţI�ܶ�S�Q㠂@ ������Y4Y�����K�L<��ۧ=��2�1`�u��Ϡ3��A�|�|8�
�4�K;��0xww�Wz
#Y8�	p��m�<]�L��K��Y�`��p����(ޒ�:��J�I߾��g��@��ק�Si�c	�n�E��\�tN�"��E�������\�Cmc�4��>�W?d��Ivk��!�t����%0_aؽ�ά����/us�����I5��Ε�X�d�f��!�c?���ֶ�e1x �T�$�f��ٝ�B+c����=\߻���vo-� &�S�f-b��ZM��~�����(������8N��m��Ǖ_��SeA�b��I�Z+5w]3����Z��B��R���_-��(��!a����A��H-���_z:�:*J�[ �a�dy\�s�v��}r`*�yd���:����Zh85�����V6�J���0��큘��hZ9Ii\i`�_�!�~8e����y��@]��r3n.1f<�jbkZH������:WG���F�zs�ՔS܇q�\,���I=�.��	ݬ�\蠖5d3°H�ߔ����/@�)�))�O�� ����������M�8F��NM�,��m��gg^��	=�)4��D��pF��\0�h'�'��hȌ?QwP��潐TR�vޑ���2ӓ��쩖�� %L@��<�YIHFN:K��lG�$2"@�ƭUJH�S|D�-E�hᩩ@��,�D�IwΡ������kF�6���H1UX����&ܻ��{ �0�U�9�ND�F����Դ��{���?4>2�?��f\,����'�ĝ�sB|��~�c\��/�2c���e�(#���v�����	D��#�l�J�ha�3��������:Gw�(G�KNL Tbh##�X���'+0KF@X@,nogC���MH(�5yjCL�T�C "����h0���}5��+�N1J�S_p��&�~�g�K4�17�R��4�����6,եo���ts�ώ�>%7�ʒ��L��c��?��R\��~�$�����֍�Z��,$�qؼ!��y��ԟ%&;����K^@�O>�c���(`^D7�4`�Q��N��h�g�=֢��@A��K+�x��N���!@�~lQ� ;��7����k��L�tM����t�8���^���4c�r�f}�!|C���N��cc��������B�a��\��k/�4���#7	�؆���<�����^��W��P��|!Դ�?<`�[RJ��N�4��E�!|�8�����S�k�tq
�� �d���U��3~���f�b�� B@�Tt|����Q�ʴ�~�}�k�W`(�{�a?Q����f�� �������i��5�tIl�§ил[�)�(�R�]VL�ȇ��*�Kre���ʐ��<�/	Bh����oX����k����G-PØ?�͑=IW�*cd����LOϯB��H��c��~RVc�?�5���ș���"y��oߕ��S1�63	/���3r��]�$��cuhS���Qd�iژ+�%�W�;�
$���z��������(�$A���Q���$��x�	_����rf����!P�j����O��$��ݟ�����![���d4�� ��p{�[J�M8��� U����
A�=�Z�T|&����_��>K󁍔S�`;Oq�b��� ��0��B̺��,H�M�X~�)CsL5�b��/E;�R����\�R�,R����2j�εl+�,0���Ir6G�hb?�1��d�Y���^�Ba��t'�8���nZ'ԃ�7��v#���!��y��^i�g�y
7QY� �*��c�k０�%�<��g�Hi��.4�W�O����Da�땈t�����
��z��������܀\�E����9��r[��J�iX���(�b�?�+,��
a,��7���("	�����3^��e�e��[�#|(�ONxZ���&!�ҁ��T������omt�"�A����J�(����?��8
��]2���ۜRN�WF��e�ޚ�+B՝Ŧ�`�i�2Az���ĊL_Ǻ����,�oh�����i��mfR�k��j�u;�/�NDd��0��H�&�_����6� T��QY+X�\���Q��l�j�ړ4�U��{�o�a���4���ɴTV�pc%qRR�Ke�����'hL@X��4��`tӐ$`��Mc�̹��kn�9�Ɲ �`ZG�yyVϷ����F-�HAD�.9�-Y��1���� 4b?�ד	��+��v�R�����*QQ9Í�J͉o���EfLG��ӛ�1��t�[�	���R��e�����<s߫-L�o�,6p���pg��D��q�ܬ?]��x��v"�2\�U"'-�=�y����m�m)�b݌����3B,�-��0{�'��7��{+�5�����i�ʺ���wi���rƺ�f���w�Q �4j!��J=��G
a�ϼĽĉ�0Ԉ�2��CkvE�2sŝ� �Gݶÿq���|y:!ʝ�75�r�Vi�ģ�c��+wC�
�JL"�-��EH�
c�<�"d���0�y���؈L����:�h����>�7<��kAT 0��4������E|�G�/άc������/�q� Ϊ>Ǣ�UW�S��B�����g��n��g6|����yqyej*���"��o3�9�b+#����[���`כ_���%�T�p��	ME��V1b�]�֑7�3���������X��
���J$ZK�H �e9<����BD�u����P��D��&�������
w�S˃(B�ʬ7�F�OHTdgBR[��`s��ڻ�Vw�Tk7�_��K��>5#1k�'�*x B��xi�k[��$���he	�.���P�!Ƽ'	W����z�iU��[#�F>�ZE`��s/��?��_���x�I�>�_�7�\�gD�l��y��7	-|ۀw���V�v)(w�����O_ q
���Z�rp�z/H|�<��P�C�t��w�@�b9d�x��:�2Cct�P�̳V���w$�zVr��@���nn��������rr*ݴ�AăK�����5!a��C��v ��}�/��`��V���,9��_��&�QO�	c����{��R\��b%�Z����O�#{O��gE${Z +�]>��_]�
p�#��u�0�F!��,�i�~z��~bX��#�^fum#es��֯�N���iW��9O�=F?V[aVB(H6�t�@S4M�fͦ1�T�YX�V �����$�1�堌����\���6+���AG�-m�o�v���+D�BG�^C��H^�s��8�:6ѐ��%By#U��|�Nl�  g�MJ�la Sr:����������T�)��(^�_
K�}��{@	�_#�:��=v }��x\+y�s��tH熿�UJ�~xNDѱ��)u�q��K �XZsZ4	[�}�1P)f|�p@���焰�&�ej���K�l�EF=��B	�&�Dߵw.�v�
%L3�A"p�y�c��f��<����ؽ�y�`��&J�B(�� ���g�k�2�����h�Y��,}	�t�޼.j��¼��Vq���42~0�J���+�6�)|��X۰����$�~6ҭ�|�{:��#��a�d�Q��cK�`�A
��6G�Eu}�T��w�+A?�A6ў��i���Ӡ�i��͕yjq���]�+|L��n�zU�;"Y�.uQ���Jd�����~,v�[���R�S�'��:��]�+��䦒�����>��N����ѱN�QM�� +X�76΃�[yϪ�ҝ܀	���'��o�?,��;��������
�V0W+���yL�u~���"�?�i���=�u1M[�s��^}���?�k���m�q�Q�'���2�r�� ����$Є��OB8R��b�]JX�k��X 9ly�@vU|Q�ˢf��2�^S���67�(�G��)�<�f�c����T����z��{�ZN�qS�?Ui�(�xO^������lκa!�i�A�o��<CZ��/���\�$�F�ͤ��LqA��5�z���H����(OI@�tD)+���̡"$֩4_�]
!1KYwh��i���.����۲��_%�}���	">?�����P���i�#�o#���������-�L��FI���w}�8n%֤�iVYz|e�x�]�I�!�@�3�Z�v�n'�J����FI}���� ��P���O�����9�x�䩃QV�ZbȺ�7��)���r2��;z \E�-���jSb�\zލ�
s.փKA��~����Y$ZY��6��	�{�Q��h����Δ�@-���:D� C�#D����"��O�:��_?N�i?gnm5���M�r�Gz�.�F��x�ۙ*��@?q�`{�`��}��U�����_��R�V����=�p-��yC|"���w7C����L��!� ,�7��A�wl@��o���b�Mpl��t+��Ů���� ��p%$X��4��wɐI�#ŷ�D�Q.�����P�Ud3�����e1*�q:փ����,ı�V��0ֈoK��t�K�IR'�g3V�s}���-7!�_��K�|-�)���D.l�ɧ�n���%J��T���K�:\7�HWQҫ��}�n!m��.�'S�1��7�3/�Lw4����%偧Ȇ�������4��T��+�f9^d���{����DY\X�����3��Ќ3�!HY]����oC�AR��
����@�+n���7僡�~�����9��q�O�16�7���y�����EJ��$���i^i�>�)>�_͟D�q�U�̳x�Y/����f��0*D�P�^v��6E/[��^1f4��
�fb3'�#p��V�;�S��c�^�-����X�0.;�ӊe� ���Cf��y�=���={�M�G��<������>�>��#�;n-H�,����)x���+��<%k);K�10Gq<#��?^@5�� �M'�)n$���%�m� EV�l�E)��A�@8-t^V�s��x%V����L�Υ��I+w(����c���*/�-�N����bt}�pTIZ���@>�D�Ƿ�a��	��>S�H	�f��b����u�pmy	��2��{�WP˿��[� �"/�:/v& m��@���� �zd^�s�(�ߊz�b>�˳,0�q�d��X�9xH� h��&v~�_��o�n){r)�NHU hT��$>�a��~�$�-���~G�a��=�B�ڙ�i�� �H�}�%�+`UPA�p����7���⠆~A������k!?y��'~J��S`�5[�.��h�1w;����Ų\�D�{���NU���H�����������dv�����"�A�ǌ¿�[C���^e�q�5>��V���	:�=k�M�|&a��%z8|S�	
>M�v����6�l=�������ʬM��2�v|%����K��&��/���"��G�u�y�&\91S�KC��ݹ�<pL�d~2�=��,ɚLI�\���n3�H�w�P�q�P�j���d�������������u���ܶ�U���y�Ը������X�`�c����.A������������X�&ʺ�����M?��Qu� 7���$�� /�5��7�=k�L�A(¡l�'\�SO!!/�Uff�PG7��6�
�X=C��
��0e�d�J4*J���v���B����X$/����-^l�ߚ�O�=g�&�$זm���I��rq0u(��"�H��&"��d����/�k���)�'D�wt���c���Y�Ӣ�
D�7�B�S�Ir|0|�n��WA��S�ݕ3��������" "%ۗ�־�Y6���/��3#D���7?��^�sǄ�l���a��I��{�����M e����e�w�o{G�8+k��P>Wls�ѣ�F�������U�e�����(5����X+��l_wGXa�Y@`%�k��~��]��5	����,�%C2*3��bXAf�&��t4��i����x��/�g��<�i�;|����k�*a����,+Tm�,�!D?���D³U}���R�S��I�l�� �l_�U�7��k�;^�X���r����
=�Ot�~�x|G.�[��p�������J=���)f�q�V�xXiM�ͼ���I�1���e��N�ϼnU �^A��%����j�j
4\���ׄ�9��!�kP�=,a`h�C��	�L�/���=�%�f]���y�	���ʇ�x��K!���qA�g��w�稧����5��z�N�����a�سx6N�9Ns�=��A,�o:�q5�H��M@S�{�6E�]��,���B���{�[I�w��x���>�"Q3˦K!��Ӎ�4��.�/V[w��tFK:���d�&�e&F�U��K��t�3e�!TU���Y��\>�>#k��CWІ%ac��6K�k�]�<M���S���G<�@`��Shdze���;�yX��H�~��ȩ�,,�A4�-�����ly+���a�(�K��� �nC%���JO��{u�\:9v�� rN=U��A����=ؕ}��eru�����;�=�Q��Ʊs[����܂J��flҲ���%"�hH쀙��T^�1j7��b՗,L�w��*iy��H�=�7��j����.�t�W��.��[�vkИ�s����!'����������a�]}�Z����:��f&s������6N!��e��� ekS�1����I��>Ԑ�����&d��=�d��Xi��Q=�L�Qɉ�O�7���Z(�I�}@H��X��0��s�$��{R�����d���	[��T����؛�k0�7�!�
�TG�Sf�2�TJ��8�&a�I~��/���zTr�{�_>�ş�j¶��9}��D���byҢ��z|zCXO/��-�O5��̙�s�2�en�qh�#�Y�q7�7g*r��� �qw�Z�-̮X�yoH��� �	RX0�X�5'-PcN��#�.��\��$��̟.3��3y��Xnfr�v�-C��jf�=u�} ��{�8���T��^喗;�c����"M;���,e���!�h��˶J;0����?�vy��
D�"�ڸ�P�u�s՗Ž��"- "�B�
ɧrHԣm����6�c��1�
`��#ܴE����1(� :������C���̏��M3>�T�,:�F�h��a�q���͢�4�P̑�:2��7)"�ykQ'&�%s�wgL���p��q\�fj�tab��cyF�ˠ��5��> �H��'h�I�!�*q��rl&y�nǡ�ꇴ@Ub��QXƱ�&!9F]kA^���ʆ �L�h�\�� q�k;��h�=�y�lWk���/q4O^\K�/�&`�3��p�eǩژ�^��uJ�U~���&8A�Q�O��	�I���pTD�c���R��w��丒��#Z�h����� �Х�F�;h,4��b�����5b>�u�{�=�?[u��uVk9'i$���ML�<U�z萴�ߦ��驟���<�%{ ��~��l�􋷐��ZA@=�	�^v�1*ߠ�]�N]�@�)�������cO�A$Ph��6����9��W��[	��uhSuѓ�a8�K�b���R�K ڠ�PI�O�ɻ� �[��j͋�����R���D*`���n��ҝ��Z1�,q�!��z;�Bݰ�OF=�x��!����ѩ�u��"���|�/���L�_NDm�B|i��	�%q�5��(�����L-u�Ce|Ŵ���	�]j� ++2�Wg�&�p���R%��5k�N��C)e����v�����H\c�pt��ԷRWd.@�y��DX$�����Q1��AV ���l2�=�����I��N~WsL�ub�mKD��v��y+̧p
���p�$��Y�P�㺌\�=��Ah�kT2�����E�S ���Cmx㳭UZ�"ˉ�:�.�Ȟ�j���RP@k���-�8l�