��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&��^L�h�m��uXҰ�O#�-�D8��})y82�E��gŞ/�,�k�F#y9�G��>m�^��N�B>P�6Ku	�Db��}�c�(�g�7�����G.ޕ�5!�����?��=���6�����A��hZL�򳬨�5DE�=v��ͨf�2,]=l�	�O\j��y%=A��y$h�P_q8�c��cF���Y�ܦ����~~m�BJ�J�sg���G�d�ul�2�P_�<@�������#�Ee��kj���J ���-����a�`;�3��Lwo��[��o:Ы��U��tET/ʭ�|�~�&��n&�acdT,C�y@������9u"��D\2KL2���t!
���' �P�pi(%,�r�"�E(�=08u��N�ld6�q}�zL�W��P�1�\���o�r�&]'��\,[Z��_�d�	VK��.Uͩ0��J�[���#ء3~ 0�c)�z_��s�
rje���M�����FI	�Zf���O@�g�ʔ�`�50��7�VP�Eȩ������B=|#G8c��9s���]5�c_����*ȹ����HtC "q�����4$<����ۊ�M��@s����Ť:����4�g
�`�!�r�Nn�\�~^��1\��6��< ��>��u���@750�Sm�ҭ���S���Jc�Ti;+2�k�Z)���ɭ5���Ώ���R��ze��M�o*�M�o�k2x�k���V�S�g�'���r��V�!+E⯓i>�WS��r_/w|��[m2�n���@-�	畑��6*< v��������	��#�j|u'pKV.|�!uXM� ƅR��6A�9p���8�p9�8!P��߭EQ�mW����4�Q%�a�za�8�o���Ț	OO��(q(��i�p�l���v��e�8�;���qS �X��kr�G�O�v�%��ؔ#q,N��fMs%��mt�$�<	�MR䗣���8�AF �s��73Xo�1��L��	݊�Ă'_�uX��V?^�{$��ih�43�/�H�`�Y�P`��� +�Xӷ(�_d_�#'5r~�t��L�+_�nKF�Gr�������:�t��C�b�ܐ+��PW�h����b�3�z?���Xn�n_4�L�VW�qM黖R3R8��ľ��{�������I�Y�(;x�/�U�?�'4�;#I2ex�����V	���@�=�BV�+�kJ�s�A\��������%:x��i�
Qɐ_L��� LS�-$W$ӗ���s�ţ2���������vkؘǪ�f�:Z���%�K�X/a�û��-��_��fx���q����;�#6H���t��sqF�T���Cjo��<صE�nn�{װi�Q�L��� 1�+���.��{�Ak��
��z��jI1&Az���ڋ�*6��I>�Q7W^D�r����>�����^��/�F����dzO~�p�hS���N���'_{�|������ϳ�ۼ3��ͮ����d��u�;O8�l�af�'���b���%>$Z0�d}����/H0q֡ c���������^�oY3ćtu��_��A��㔄�����}�p��{0*�!�)��K��%������y��B��;�ձK#'|���C���HD�P@�ֿ��~�y�XϷ~'Z�f�����(2�%z���Sʥ���������95����W�כ"x��v�Z��#�2ݓvy#Z��R��2hTp8������]MX[�əTY��L���Ȯ"��Yu�*�ՙ��9�cNe"(�Tn_����S�G�E��૳sp�$PS\1d��&�-`?�@y�<�2��]}�&Bt�l��?��o�Z�蠃a�w��T��ɇ�yvp.j���춽^u�[j�fU��S0��BY~�A���󤊬��+���=��c�6ͣkEH0[�!���,�d�c�g��R�
�{�){D�C�HjGk����d�L� ZM���c��Ö�gD�$�_�ܗ�N�
�
Ϥ��&f��IE��p4�B��:�BXN�˳��>^�����`�`͎���i� ����L�MA
&tR�|�`
���^z��I�����?t�Ӊw��m �,�\�θ�v���ӿ�8�I�8�8^t.:��n�:2:��e.�̓C>�����3�F�#�w(D�5maAL ja�?)7���pk�q,���y+�����z�K�5�\�[B�"v�ǧ}�2/q87>/*Z��WtXtj#?�c'� ��ñ�WGCF>v����E�`��{0�~�S�m���t�BR�����nt��V����?R�Ȁ!Ysֆ�x����cٿk��)bR�"x��E�4��w���3���q�jj����w�X��rH�Y�I�X�|i~b\��ef�:ʜB�)���X�i�ƁfU���<�z�%����!�p�w�0��.�i�E�)�n+K7)���BA��[�x�L�	F�f��f@�-�YO��o1��߉|�S�N�H7���_�a�oHN�U��|676��;��EV��\m߬��;'G;r*�)I�Lg�͔�V��tD8�)��*��w�Iu��}�:�ӡ�C��"�rc�����ֆ��,cT�*Y:.#?�P=�9s�	;������%c,��,H�)q\�ȵr���Ȱ�,!��	���l"d��Gb(]�dm)$�s� �N�z~�3J�F���HOD�s��4�����^}��S^㐖�����X��3��E�:��.�w�BKi�Va��7�|a�
��ړ�6M��a>J�屐�ȇA���g�)

��b��<��#<g������M�P�j����-H>~�h�*-�V��$���B��?
LC9̉=�m�?����(_q8�l�7������>�����(y��7�}����_����T�9u?ك�1K���� �;l��\܃�����I|���4�uD�8Oԍ�v�P8g]R?:�o/aNGI��[��f�o�۾�tR ���tխ�8e-*�q=w� ��fR�\�ɛ�<���o�cF��d�u�֐��W$�-�cX��+�'&�T�H�L&B�.�.Š�����e��i�����Y�����Klt]�N����>��i�AԜ��pQBv��'���:�vD']�>bM��v�uM�S`\���@�޻T��=[5的7�-z;�6��n}��@U�,i�+��@���.o���T}=i-���<���Z�{�p� �>�W��Sy�����h%N�e+��,TbӠ4y]�����<ξլ9����h�eꙦ_�\�veF�=�>�4Y0,h�V��ԁ�hi���AX��}���K��-�y��{Йl��NB��I)�k6���K������ɴ�ջL�p̯y8�����v8��z�]z�j?q��c/�!��}�v���7v}P%u��>�iq��t�G3�⤷�7�ÖV�Ĭ�?��"��/XR[��zz"{W�^���M
�"AKq�/^����LGҶ�Z��p���G�4������r�[�P���ϻؠm���7o���>7�k��p���6ds���&�u��5�P&��7p$<
�J/��v�����Q�/c��e���F�o����G^?�c9$�J����\���Ɵ�`ޤ8�D��$�N���o�@C*��2R^^����Kz��m����/R�(n�Β����x�L�	ԅ��+��W� v���1ǪU�˩#}�#��/�_}�T�"|	������uE�ADj�����o�����XXR:
��R�u�.a�P��6��x�:�Tk��4����P�����^���n[i!�A�y���e��U�u�Zm|��&t&��l���Я�*�da}�n��3��	T�/�,�7����-��#3S�� $��E�Pl<���k�2�<�P¸��fIkc�:p#b����<�����=�#s�?�F���-�<���M�P`�c�jv_�3bnH*���Ň��@Ƞ!a!@ܣ�o�4WO�bu{V�Z��EM<�Ef�y��C��� �#��^j��bR��ZqQs;�J���B�R�����B�N��v�D���ֆ��S�u$���X�:vY���GQ������L�����f�En��X�F��'�q�H��$�vƓ~�Y�|�9��ڎM(����_)���~
W���?�0��>��!�!������K��h�N�6{�dd��>b�A���!O|�Jlq!ʃ�U�D&;S�Ɋ��zߑ�C8K�����犀�,V�Ă^�g�5��,;�hA�㪾�v`�w�r%*U��׉?�-0m�q��������n��Zr��_�*� R�n���X.���G�MX�bB�~)�S{P@*K�XI�$*���؆��c����&:�?���k��>���jC�_=���S`��[�焑�-o�E?�U� �W&��Kd�e2NFͦ��Jy�hQa~L���"i��,�0n~�T4h]{���'��7Cb�H�u�x1�YӨn&������^l�2q������Xve�%b�����u
�
;z����Ճ�2���2w�؟����"��~N�-�e�:�TOp�H���;5*X �rѫ�W4��G�-U=2	/Fˤw�D���Hz�%�..�����^ͯo!��C*VɀG�}n���Z�#�'��4>R��0��>0t�w+���ھ'�}d��<��5	��rs���w1�O�?�h�!����XN>�s��̯��It:f�O�e_ �f�K+^�(s��a7>�,LΑ}C�bV◑i���{4���VH�!r��Q�Ɂ��(k�{�����~�*0��ʆ���f�9ی��p7'3՜�C?��� ��?��c@���İ{���od)��';ɪ'qk��0Wz!S`�� ?�`���e�l\}��P�R b��mj�fO�F�����=lfh���ѻI���l��V��Ph���~���Ҵ27;:GMf���F�N��c>�0��F��p�������2�o6�|���>G(ȏ�-�܉��/	T9����0�$����<�`m�z0��F� �!��N�����I\"��j�ח*�etG �o\��d	�\�<($�TSk�˕'Q��{ոFj��5d1�����C�l�2�*���?/�
h���'�$��HwZ�F���%�O?34������1�K�R���W��\��
��ݛf��4`3�0D�m�� �6NzP�&����)&;C� ]ۦ�x�{ə�
z�>0t�����y��kw���I0Ҁ��O��T�(���iଋ@��48�I�^eh�j�-�,��fv�M�>�?<p�J���珖�Or�s�4Ȇ5����+�D4s35��k�IX�p���]g�*`�C����~�>��k51�~�Uq@]������-�DҰL�#X�o~�&�%ǳX�F���F���v�V����u&ҁ��w�H�,�h��� �Q�&�{<��J��uWer�Y�_b��U�XsF���a�`��y��������L�ּDlj��l�����G<Z�N�U ����D�\��yWi'�:��<5�fR�;̥ŝk���i�-�����7sp[i�IЇ�ʓ��X�����<�c2 2�������Ze�%|�ta^$=F�A�G�G �� z8p�a[Jir�\�6�ۺ�9��Ę/&_�_ �%U��'Ks�_��f��֭]��]JOE�-Ma����؈�-��]X��>���O7yh��K<�7P;��WN��{����u&�C��W�E�b��}-r !�C)6Μ�qU�����UF��J+z�nr"����Bc<�k	�p�wn ��gw/OmˎxY���|��B������]�?����,|��
�yVP�E*��1�[@������N=�k���x��^RD�(Rt_����D��_�:��ҙ��3h�4�p=����c*�����K*�J�u��]�T�y�W�p����q�>L���̆+��B�8��n������B�8|�/���wC��4T��Y�H�r�����y�z�4i:ud)'��|����~�)�����>��۸ְ�?!�>���U�����QJ��-N>���(�:V�#s��<G��W�����Ѓ��f��Hp��h;��J{����^�i�r0C�F	�;8n�W7�Ԟ����J�+����ovޱ�26��OX1��Ϫ W������a��= �f�,k���`"�qhA��M�ǐ����\�O�x�͏�BXG�`�%K��jꠗ�߈��5 ��}�\l��������Spn�xՉv�˲%��qe�C��j�$͔�����c�&a��Pw���8w5(
�򗫺�X5�Y�,4i�u��8�k��:O]�6Wra�a%��h��RI)mv�i1qbeF%9f\6 ;�u�Z��e�1ɺ}�>d�ui_�j"��.��Op{��z�s)	`�b��)]�� �"�'�fi:ov�NЦsw���`�fUr��~�Dgq���y�v�ڗj��뢻G�W9���̓�[��k��6��!���x1�m!��W��mG<J����H����w{0���!� ��{ט��@�97T��E�)�aiO+�#��2�̤�հ��i�7�ǰS�*5o���P(JM�'?p���q��`�_v�c)̦�J�,
(�},H�S��F�f:�MK5MU��E(-�@�ؤ4�,(N��S�ɼ#�F�tF�	�ʈ����;�~sŦ,��΀��)Pcpـ9�mN����_��'�y�P�Ƙ���a��/��^�7��;�ߦ>�{��J)#�� ��r{d�靓j��G������k��l~��Yդm���AqJ�,�?WD�vz�`��@�-V
���rtA�����p4�7�I<�Y
i5n�Vn0��b��ڱ�f�!h��I��9<���?Ƣ��Qs1����-���}�r��#:���q:փ�WcH~�R�B����(��^Z��޲�T���m>H,��ʦ�M8��!n~5�C�)`'�6 ���Pϊ8��b��z���LS���:x�n�M=H��떼��(CJ�5m�����A��!NSҹ��7�0�h\,���h� ��sI�Q����Gb�|�DSL˴�bR2qѤ�̪k3O��!>H���3+��È�&)A�n���zIj���k�cX�că���_6�����%"������a��	�B���	cg�7��������a���"�=Vƶly��l]�p�]�x�)�U��q�6Og�Cф�'���-5�q��U�7���b}��槰}�ڤT��w��*�v�e��)�)%}q���H�k��|hoa�����J�[vDZ^���m�M�^p����C�)i@_�����gl4��1��Y?|%��c�Qu:�7�q�|�ɹ�b�yAr۬�b�[���tۮO|ft�"4�BA�u�珂���0��
���N�����/[��#�{�N�c�-k�慯C�8�HI���M����ix���� �}T��@��A�WWFV9q�	�y@W��֋ɿV�`���r��(v�i*:82�ŕ3�7�B�O����c���?$�|S���-���3��dJ������ܔ?��/�&n�"�*JˎA@�v�ĸ�1j�"t��m�[�Q�u7_�p�ng��)�w����l8!G����m���4�H� �r|��y�)w{ͺU���+H�SFD�0<���e�zê�T�_��Q�[k.��7����T����D�ǵ�[�_�����:eyC-c��P-Y����������FX{����ҏ�	�.[n�Ꮋ���d��a:xc�:z�Ax4��w�?�+'�b(�H��I�k̥�f�}9ҙ���tvrG�w�וPS].@���,�������ޢ<f�bL�u4������±��ϻ-?�-�ꨔ�{8���|��=���nN�?����E!UzA�x�HҰ�>�6B�:�3��t���
�3p�l�P�M�����	�j�n�J�I�=�SR�җ[��H�&����u)�ғ��F�,��α��[��)���I;Q	���5C�5�0A
"uzn�"g�_��qZz^���y8��|K�`���W�{�p��@҇�;�q]�YN~]%iqYe���Avaeh�Lh"���Q�hړlq�S��2cc�ލ��{U�$�2��n��wAIa��7Y�Ps	H���!�l���E#xAA��AuhS���^7)���I����UE��.2�N);�֧�����̀�Jw á�
�caEQ_�.�=�5�e%���qx�WD�@���K�\Ĭ�6��RN� {�h�VQ;|�{���| X��H�|9=��f�p��C�O ![aY1��1=pW=d�N����9��m.�uqD����R�/�2x5�~�~^10h	�w\����I :\���Ѐ0��Y!��[F2��P����)����R�NF����u�Q�2X^o����lB�g���=ջ�^�X��dR�/}@9�F���)H��F�*>�,� o6��̅���Α����4�H"\O���l��F�p���g�}�����BOo*97!N�z2�4	(N��2��X�)�[�д����s�
�aQc�מd��aָB��KQ�!�~� [R��UFF
��n��5ؠE����UP�+�Y%O��g� ����ӳ�e�^�g�3`������m��ǯ#���g��� I�	�YY٠,��=㭠�H�.�n�s�%z��#����l�M5�v��"ͩ��dzŗ)���Kh�Dc_m�M:!'"��[$w�`5�����O�GMZv�@���f؞Y�ǩ
������?n�L���e����T5����;�f�\�ɷ�i�T�㞛p���M
������	��7�1�'y'OA���U�z��	�?J%<�e��2���p�fا��V�g�iJ}��"?�D����C&m/��������	��qX|�q�o��Q�|�#�����+%�����ETE�\�_���R�Mz�;�`1{��Pӷ���ڨ-er&Mk2b��kV�U8�6���E�|,`l�|}!���֮�f�|-rƆߗs�Ŋ���4����ɔ�Y9���/��Dej>�޲õ���a��Tn�xz�R&�^E��	���������\�S��V��巓4�q ڲ�\���4����ە{����f��ra����.����J̺�3��,{Se��Ź����A&]��qj�WF�5*��-��&�$�uv롁��:j��R��*\��e����s,>H;�-��}�������N�M�6y�`gcjW�B ��]Pe<i9/y�;Ǚz�+�++��eOa�z^	����AAR�h�8]�����\�A���Rw�i؇�'��v��5+[�c8}�	.��g�=�M7�:Sу2���$����'R:�Yx�ı1 ��?�ɥt�#�h�؍H��=�&�/sY�'�F���e�n��v�U�9�P��R��8uE�X
��==���Zf�:�D�·[dB̳�sQb��6��.�~m���+�Eʡ�)��a:��	��~��N%S�z�>�f�>Q �~P$o�z�R��_�e�p�[��n��i�ː0��r��eW�PO��_���C�+A'+�Egt�*G�y68�^�ԈTpi]��uW�٪@�F��yJ����an�ސ[<DW�Y��Mn l���#��k�[�o���L�U32���H�l�ꔔjCӉ�8G�CiYf���K'#��{�:�7V�[�=e���K?����B�<dy/�7r��t�3��q�?���J�s�ENs�cGPZ���W*(<��IXL�Zɩ��:�d�#ҽ~�'�Cc�U�Lp�+����v�����]��[��Z4`�p�Z;�[I%enU��p�`��'K��v�U���_�з��5�$5ϋ!�ڎ��ۤ���9���O��R���e�70iRΥ9�,w4+@��ڎAȝ#f���o�6���3QI�͈�^g�\���͏m-�%q�Mnb�sm��9�����f�V������H���|"iqr$,јt_�Į�L46[� ��;�heϺ��NH�#s��g�2v8Ѣ�H
ܕHcx�SH]Y�t�n����1��0�x�?�JF��ɘ�R�}���[,�ޕ\%��*��=�Vy�}dU���@s���8�?
Y�w���C�
(��̌�7+�$��U1�>S;Ƨ�Аׁ^Ό�rI�n�i�k[S'�Cpybf�5��ma��z4+�+D[Ă\S�=�*��z�X��kWOI�7�B�A~P�"����T��S��c�2��+#U��6N߂�v���;9�q�B�E+�$�<.��p�U4�͆�9d�qi�-� ��[ԛ�̧�d8\2���/S�8  �xz���YM�B�Eu��D���t;���hi��J�z��j:�p��� <Ӗh�����K^jb+��Q��m�����#����ƝYl��8*[�˴Hb�N�������E=d\���<`�w��I�L�K���r����<��	�w5,�O^鑆���?�lf��`��^ǔTӲ��:ф����'8t*�|P_�$�ަ�����t-�+��|��S�� ��ޏ	�<3'���h�;'RcO�)����̔����W��E�|uJ� �_d�#�]�/��0�:UגnC.�A����/M^B��wd��˶���i��MGǖ�������sw������S�]3;�w�'3����;�5򓸺B��kZz�99�x8A\�_,���"1�c��g�6�еtiR��C,�IX?�����5��bP	�'�Ȏ#=�����p؜ڮZx?ҡ�=k�����2WU�f��k���b�B��5���G�
�|���(�k��c�'qT3��`���6��x�I:v� ���%>�*��¢��K��VZǚ��/�C9�L��v���2��=xR8R��s��n���.��7ڳzɸ�A$��i+��`��y�p P�j��NLy�.; ����h�
y�T���bk��ud�wa�*��h6"��X2+yX��Ӛ5ƕ�V_k1��fWt�s��9iI����Q�4���(�7D�ː�j$��#Yx���pބ�!��%�_f�xs3�"s�|o����ߒ,]�
�S��͗Nl{�")A=%�,e�z���(f�o�����x%��=le�6C�z����Ua������.� Nû8M�>���iV�G
�k�`�p0E�����;kƇ�;��<o*Q���_�)��k��ŀ�\���$q��\��+��8�+�-��ړ��6|��'�\�'V��h���1W���*JE������4<	����I
ٯ��{����{�;N�.-2dYGۿ:���m�
;#�WÈw�����!�&�T<��{i��G���W��&�^Ny?�?�:���,�g����~��[ԩݲ�44�p7j��)��P��Sg����z���Z��;Q/���R�r���А�If�}�q\{6��$�Z\���E񧑨�Ʀ~�����_kmYT@�n���JI���~]7l��[�7n�2�_��oYY���L��ʆϞ28������K�E�[��tog�[�,��϶�1_�)�*S�$	J�ޗ���LW�ʺ��ar���\�e4�`*pa~�)�4-=�P:f�:�@7�A�h(��o�*��Ű��=P���f�W��S*�`�NG�.1��E�"5"��p|+¹ ��$l^�#���Q�7|�$�y�b�;��f5�wi�-�j�B����2m�Axjb�2�W��-���C^�T��δ�W�Z��p֊�Z,W'���k���x�7�~ž�,�K�(���q,���\�E�/]w6)yPr�̱0O�#�����r���E[�1��B^e;�nx���#m5mn�/�۬Y�����%I�鍷�Yo�^�1��B6\T��y9/v=ZiB��6�Fg�˵����h����A�5ɩ6��`l~+��k�K�ɖrt+/zLmz��a�d/��~�#;b	�ݮ ӝ��_���~]�V�1� �{����,����󫔺������L�\V걥����et��?(1�D�Z8:c;��Ŋ�ݧ��O?ϋ����6۬ˬUX���qm���C#�eW{���/ݐ.�(�p���{ʶ��Oqg����h��P<hT0d�!mdVڏ��Z�P!�te�N_2�^\����l�+?�?%�$I�;h�c�G�NN�~4�$�{�ÁU}b��`d�2���S�!]�ൗTP��%��l�[�	�X��4ӡ�)U�̈�v�D�!���i��9��n�5�>���
���Z�B��d�.|9�ՐlE�2C gF�����ۯ8�;!�����$�f7<OwW+��/�=|kpAW�Q/VZ-r&T���k��6\8:�ۦ&#�V��04\�J�7xp���~�_{H�:Y�EeS����IԆ����$fsbg���FI�mb�x��U4<�5)*,˛q����\�c�+�3|p��3RRz�Z#A�SK��C�K-�?���Ā�T5U��5���	�@�`�|9k+�"�]/Li���}&�G8��R�ӓ�I�ڢH=�� d���x[��χ��_yI_XK~rcR9���	yn`N�8(��
�r��o��nu&��%%��u��eo�����'r1�)Q�N��-|��B/�V�M7�t�V,�X��ز��<i~V��@p���'�X��g6�c��ї�%�������BtV���l�D\'�r����Tl�m`�![Y)��d��@j�xY6�fۍO�nҜ^8H8�?�R��q�T�.���)v��s�%~bj!�i5���%��r�	`T�Pj�Y.O�D}�`GU>a����G4�4��7��L�Gln�֙BY�5��Ez�5�p֔~x�Z���?�w1�m�V�*����T����W�0ɲ��F�8�v(<����Na���1���0���_H��-������t��-�zV}�0C�NZ�M�ew��D��yj�k�&��d{`�s�A8��+�Zf<E��� HsZ���"�L<��03�y�#�5��c�\2#0��AD)3���wj�K=N�X��f�Z�6����Ԇ+�.U;H%�-���l��/��p�}&�;}�/�[pD�ă�� &r�\��F�����j�)�H�-cH2�=����:C>�	���(k�}uT٥
����h+凉8�j��܃?jTt�	�x�%u6b�鐢]H����4lM,4kn8�ʌ6%����`&��L@G+���Ѩ����]���YZO��_}l)"_���3Be�����Rc�k���2�BC�߄/4Ft�@�����R����N��i:� *�7�w8(F��� "y&ւ������F��U�ɯ5 ��-A'�`QAPZP��`k�߀��}�<��)�枙����9�R[4= =�`1kh��|!���RF�j�z�m��T*z�S��>o�����ܕB�A���f�ɧ�sU�؋y��Bo���n�ޯj��xO�71ߤ�t�WP�'���tK��jާ��7�S����G��P����%���*���̚�8I=eؽ�X"��b4��/�3LP/$y{�I@^����p��Re��v�����bFhz�D��v_c��-"���l,�݆yl�B��,<ƯP��TDN�ddY�:��]�E7��N��`	«��2��O�����7�@F�k� ���p��jM�=*�0v}���[�ۓ]^�u7�+e��k�^�����k�F�]��� ~#����Aۆ�N���}߈Vo��z[�#h.v?����7��1�������x ��U&���"�G���X��:X�8��ؘ�e���s��f�!�<7_!��C�\�6�2�{˥hy*�8_N���y�lU#Yn�eǳǝ�ϡ8o�̄�x��i^8���1	����Th4���>�<&K�-+sH��_�'��c쿦i��e��<�r
+}D`GU�~��>tR����i6�c=�8�N��| tz���Ӟ'�q����߂X����$FE��'EX��?����w�"�0��\o�{�+�J'-�W��GǸ������N�x�49-�x�����`����U���xíV�*��D�V&�\8�q�kФ��'�����>z�	�6>QW�?���q���[WFM	7f@}�vOy�� *�	c�.��b�w�cW�+�)��"mo&,u������a��;f\U3b.*�{r�~�|rh嬎�i��}�`n��&��rt)��B�x�S9FF��6M$�f�yI5s7�d������l�c�J��'��"�������^�2��>8m���L�o��Uz]��qZ]Rd4�����׶P,wX��n��uD�N�_�z�34o��F۷����z��|k�"�Ϩ\�^r���/���J�{��l�
��������Ӌ;�]��U�j�:_����$�w����Gəɉ�G=Ag��EO�Tj�$u1!�/����I�)^`����UW�F�C�ȑ�EP�:���0�8�a�����&�@2�Q��C����q��P�&�4k�s��i�r(�HR=L�M��;����6g���\ �'���;p�h �k�h@�9���M�i�n_���!�g�[�ib[]���B�Z����1
T�}��]	`�%�z�иÏ��dp��b}�Wd���#��v�rr�#}�՚Q7��o�;�n{�/�ʗS���f���6�H������Ct+2!Q��{������/5:A
��#���=�s���k`y�̓*~O��e�ǰ?T���p��O�6b��Z���^�{�S#=��}����\,�Y���_�̓zUmD�S��^\xkn#��\W����P"�0�HS2l>t����ށh�=]70U��rVY�����V+?/������dpH~�&﹜����BsӯB��r�ZF쮻cb��|j�Ȯ���}�߻^R`�Ή��zT}��m}�W�q%F���T�H� U �fϢcF�Ph�#DD�o���-�FV�#oWl ��7F5��vWR�DE�%"��nD�e��j!�nrH�q��$�#z
(}�-����F�~E2��g�'�� ��{<OAW��<Q�Ư,/��8��Z��0[O-��R��Z<Y�8*�F�c'+�]���+z�k7P�nF���B�W���%`��	���������O?Bڱ��>8�7��z�3��~60�6���E㘦�h�����Y��~���t� �ɪ�����鎪}R��?Hm�Uƾ�|��ַݧ���X�h핶�Z(y�����ZN�?�Y����B������zۑ}�7���=�
U,����R?��7K����؅Ȃ1о��p��K�B�����:�S�՟�� �r���E�C�G���a�� 	qԎ�O��'�D�!Ӑ��"�j4&��.gG����X%]����~G�Rͫؗ/��;WA���j(�"��#�\�����]�}�P��)��,�a�>�˸��C�VV�VH�=�.���}��vJ���7\;aGo���.C��.�X�������}I���pE��Z~�Ru"�wv��S�q��5�4���I٭im��y@H1���zX����~�S+�s������FeyMWt�89��ucs�G��/�])����l�S�2�x���~?Q�kuH���m~�a(\i���%�S���_~D��������k%{rB����Ѐ����?�����֘s�'1�DB�<�g��U�KdGg��WI��~袲Oڤ�>�fO��:��T'��D�(7J8.ъ :T����D;K���<X�۵���f��vo��T�a�T��*S<7Y�M���������/��c�,&)��gk1b���$��͉���;��ˉ�Ϩl�5$��t�l����c��$�H��0TRhq����Z��I�RG��7��҈w�ht1��Ok���J�
O��$��f�mU����M���8�|���zoT��y���s�?�kI��#[�]��������i��!p4�,w�r��_��K��O��/-������%s���q��j%V'61�� KnV'�]1���6�n�Ѣ� �i-�8J8�Z� �����I̿�{�{��R �Eo�2Yy�E�kBr]qp�g�3S^��?����,���$<��!�bz�<7L�4	@�� G��z��9�"�^�,��镕Ȧ�(K��[Y�*�.K�`��Oz�t�0��S�1��)� ���;:p��A,@ �e�����-��
c?|D�}�B�i�-r�R*y<g��E�	.�j0���ą�����WN��'��������A�st#a�{���
����/�ɬCWbv�JÁ���S�7�� >�z�*�?/��d�Z��+�蜇i�I��gP����*m��s�*V�B��/ibb��M��[T���m������N�x�N��ؠ�<�z���>~F�*�b�m�����YR���۸ޔ�G�犞 �;T�'Ħ�����_/{�����	I��q��������+pgzHa��h��9����h��F��"��mU։O�#y�FJ[|Tٝ�3g��w[c�7b`_H�Pj11�|xg@]�' }ܘ���u�3�b��}W��[ok78�;UoN\�s�`���D�Wɉ�	���MĄ/����N��D��%v�
v��v�k�sq�WRK�56?r���J�k�_2
춎�ܹ%l�6���;^bx���(����"���dn÷&W�1`c��
?bY��g�]���H�%��@T��dp���\�����/V��^m���*�g��N%4����N�1uR&�Q�R��)N�wzu�%�'�!	�=Y�lP��aQ
 ��I��e�t*��F`V�ܶ�v)��;�9u�xFoa��^�����ȿx'��߿�`��`�٣�6�G緷��	�;;�37��U�\K�f��
W)����(��h����O��'�[2�n:�M�ȕڃ?�*+t���c ��ǯ��k�W�\\RH$�7��#M��n��?b�|pW��jC��?\_k�3�G9�*4iE���8T�����8v�v�:�J-��b4��J�R��� .���(��}q4Z�MK,��̈���B� ��g�#��6"��(Ob̝_;~��e���%ѴR�T�R�%��B*��O%J���Bx[2+�ޤ��R��K�?hKg!SȸCJ�jx�l�k0oH�Y??�{m+T/Z����v����!vY�؟b�R3lHX�� �39B�wOQ5v�%?cF�M ő� k[T,��2#�Mw)�Q|WN�cv��r�rM�_MՉ�i"���J�9�R?���]�<�Ǩ��2j�:��A-�)������M#�CcmJ�a�@;Pt]�~����,;�)v���4�w���b�9 K�����4{\�&� n)�Fȷ�y�OZ��&FϝE�X1_.�=���)%��q�&?��s�(?���n%�� @�ɜ����z�	���2#I��K���.��س|J~�_��,F�0>���Hɉ� ���z�r���qʝ�|S�S#�������Œ�pS��O�������tlbuX��A��|���~�+P����Hܛh|`�ӖE�N�]��v��I���@���m�e��C^�,�J�6Õ��+������Оk<c�SH�ƭJQ0�%k
�������ꅹ��Bׂ�ߵ�_~�������A٪�]�?8�X��E����cm�����&j�|�Y!Ƥ�"`_����^UAT�;�㕖����8�Z�����9�4�,'�I���^��������������|%������ނ�qY�E��R���� p���`WXnJ HQ�Z�� *4 ��� �x�с)��>���Y��\Z]�:BT����0��i?Y�������z{�B� <sK�����k5XѢ~��#H�u�.	l�w��`Y|�x��>���%����e&�r�(j��x^kf���vh"���a����x�@/�7-�N;FXG_{iW/��>��o�-	�;�k>D�q�DGz�j�����b)����8s"�V�&��ge�D�g�]RwjZ���MFv�m&L#�4\-Ъꂏ�"Z i�ē:QE���^D{c������t��m��X�$�]���wgn:v)�RKU+�'�A�wʃ�7:�@���{���MKQ�r��.(�����iq�o����e\KJ����}��uԲ䉓p��\�AP}/��2�`B��Q��$��������� ���ɇ]+��'�����g�nk��]�&h�k�SmC~���;���C�+.tY�Q���u�����*����nEU�_�6����ۨV �;?���Y�$ �P�����kiмV!�wR1��U)��w���ƨ�I�5�N%�`�sZ����<����c�n�z"��TF�!�̪_]�:�PSQZ�q{To��V҇��zr5ծ��}V �9aR��Q�ǧl��oJ3�Ŭ��jT��2����qטVr��g����gs��2s�m�߳��ӳj�fa�]��&���-T�bc!�Rd;�4�#��y�[��M_UeL e���t���*��>ae!� g�n�4��a�F��/_�+��3��z�ۏ^��F�.CK�bR'c��b�����b�������DZ�J���{b:Y�
�&ɏ���n�>��d���G��s�m0Z{ڪ��SJ��1آwTP�
G�>���J��A�>:��^�3m���v����prKk���Mft����ދ��$G�'�X���d����V3i����*���Y"�d��v���,F@������r�c�����s���
Ѐ�uW�LGO!bU.�3�b2�,�S����3@g��{����\)LR�aT�8�>�J��%����)`������^�����h�\@S�k�t�}�6�&�Mb�ӹ��]�^WR��}�_�ϋ+��.�+2sH��y��e�K@����!N�J� �v<�9�u��_.P��&��w`����=M�Z�FI`�Ҙh+Y;Z'�P4c(=�bsړ�e>��i�@.z�ϛԈ�k�T�!��AC�塊��+2�#;Fyr�K}Y$GV����͕�������/�}����9��,�0��9<���o)���b��=��i �L�E�C�'r)Y"��ɟ-�"�s���nʄ�A��� ��u�F�o7�`%˗����^��0��b�B/� T���)�&����rn�[^����k|&�I��`���꺕�8��q�ss��,6HX��wZ�9k��+�4U%M6�_.��{��>�e�K��?�-���ǭ�_��V��`��o�+$�0757���i�3����L�*\.�M&Hze��Ǡ����yX�̼/�U4{/�6v�=	�7�� �����H�d��_t�m���oc�^�߳+�]�
R/Ѷ,�'���6;�-��!z�ux�Fh*��$1 ��A`#��V&�VT�P*�?��pœ�DM�@�kt�݉]�Wo��Jɨ�"?���)�Da�X��Ʒhf�k:��4u<W�/;�����&BD��1�m�5�􄹞���w�
�!��[� ckuZaL�Tx�B�{%��I�ӻJ��^z�!o`}��R�٣�3����:��/[N$�BD�&�ϡ:z�@a�s�M�� N�T+�0c
��V)&���w�=*�f4݉ξ�l���"�RH�<��ce�z�W�-�lG{T.���~M&0+Z��r]u��"Ƽ��Q�Jøꮲ��yPƨ$��7�k�S���Jo1H�]�κ�ʪj�ߌ�EQ��/�*�}MHk#V^�8#��Y��i�޿~Sj��!��E��)N�1�_|��bd� �����Z�u��f�o�y�Y�,[�6:}��ꮏ����4v%"2�w����=,�'�ē��6eJe�j����ǣ*�Jf���~��O�Fڞ&�����TI,E�|t5�S�/U�Z���@\���#��+����P��=D&b��m�Y:�Y��lj��dyC�G&+lHM�=XM�<�0�l�K��G�����~���qXr�"��g춤D^,<�Q�[=gI���%x����eN&-wX�b��_���d�~A�W��4��+�_���Zh~ ��v�A(K����,��\v¤�<��1��8P-Ƥ��$�s�Mr����W��VRn�f�}]�һ��
�~	>]������M���3\��ehb��ͨ=���F<ZF;��
F&�·g�M�r1~��<�M��A�ܐ� ;Y%�:R�/h�l����i��.KD7�O�p�F�GKc")�X���Pö��+ �H�& ���oX�(��l��H)`��^�����k���p>l>���8O��D�ӣ�,����eQ���I�X�<;�n��\��c�x��3��v'^E�T�����Bև�4�b���{zk�Y�aX�Wx�B��H{��� wa� !��A96Y�w��$�T<'�L�#���'�8���t��ֳ����(!97[ �0�ї��{�Z��_�c�Ѯ�340��~��Q��\�b��7�o
x�,?>�R�׶A`��#���%ӑ��!�H��nH|�FtZg���.p/I���ϋ��݌W������n�^�18��#��K��|��'��lT�b]T=�4�L�jT*�����s�3R3�f$/������V�̇�&0�C���zy3:ͳf��l�{<wv�s
na�sg�!��#i^���M$�|��7��I�I�^�V�6ࡶ-DiI��AH�_ݿ�8&)A�O�$>���`[�v�����60�$m&nL^�����#h��IA�i�Ql@u?A�����F/z��@��Ãa���M�q��`:�Ipm�֬#*����6��0�)Z�Ҙİ�h�FY�ljO�\x����ء��Za��P���P�ѹYt��0zu]��c9�X��{�EF�t;�����ϭ�������,{�EC���]-Rl������P
s=�x-\f$%Vx|V�<����]מ'�����/��B�%�.�5�Zt�d�4���v��F��e<APs�IG�\ ��5��鈣�V��c8!t����ШOq�8��j��7����Ce� �l[k����A����0�`���8��d�-��e��j}���r�Qء��CWS%�c��9,�����z������/':�g ^ς6�śd�ڟ%4�F}M�8L|�p�J�&���|ыE��V�|xB�EY�[��YC�-��)��b���W+�ϥŢ�J'�c�c���^ePW$��O8�(q�t�����À�?�!仺�~�$��R.� �fDXIk,x����h�}�	�0r$^��W�=�4������LKp�����+)�����uK:4���q�$�Z�.F��bxjl�hb��.J=��8Ⱥc���}8�S.N��h�Qe"��I)a=���(����d�b�G���q`���#h��͇ ��z��:�o�$���I�*4�����F��� ���~��>>;��|�j��R8<<�Ͽ��d[&?�o�1�RQ���j.�.fث�!z�>������b�F[��e�r&�u�����ԁXr����6��ʹ���Ve9O��,�vh0abKD?$��m�r�4��ɪBv� �
 �#��;���U�E}]��=	���?��U>�ϒʇp@D�(�y�����Q�s�}\��7�[?B��?G��,y���I"ߝ¤���}H�HP1՜nY#�X��y9 ��HH�W ����CH�d�+y3�j��;ĕ����Br����wb�����'RhI/D��T)���29�8�}|L����Z5�s���Ȑ]��W|�Wd]�5��V3=v�L�
R�ZT|k=��~��tV.���o���Y��x�[�	������� t�'3��{��V����Ң&*e���
 �V�i-�}�ǆ�����Sm��n�`b����!�����R�JZe���*�A��񋉟�o�Ͱ{�v��Y��]��s~�;��K��(Qs ��גaO3j��vVA�ڥh���p�Y�".�r�1�#5R]�&&�6h]�}ǗD�
���1<s��Й+r�J�\��jH�
>m����l�|��'�ؓ��kR>Q�1}������wt'��8,���%�U���H]EZ�oV����í�y9���;,��
��hы\7�6�Q���@b�[-W�ʕ8��Z��"l��X�\{<c��;u�6c�M��.=���0��YfR6��z'%U��N�ъ	����#^�
i�a�4^�-D��e03P�GY{~G)U�oD忓`+���x�Xk;i��/�*̅ު�L%!�Lz�:(��b�v7����j͠B����y���?�_��	g�9�5���Bq�~,�ITꀡ�hrhǩ.����F����<W? v�vXs���J��fo�n���#j\r��u��۱	ݺ�Һ��Ӡ >GCs�G�:�/w�m�c����o{@"�ğ��V"$͗�]�hw%��/��X�b��	��uuAҪ!:X	�����l��u���|�bD����"����R�v��_t��ZΎ{79-��Ć��#�2NXq/��_M��4���p[{���Z�=�@Jq��f&t�� ��(�� �s��"_���˶�:/-�j��9�τ]�sa!ĸwe�J=/ER~u�XW�5��ϣ,�̑*������CP�أ�$����A�{���F��J� (,vɯ��GÚFp�/��S^J�bD-Ж֝��1\�C�`e��Ά�iK4�m��K.�F��_׺*.zR];��M��ݤ*<Fm��R>�0���Ꚋ4�N=��B4H=�a�_3i(HjA������)�5��~}F�\�-�l�V�~��d�]Q�̷�M��!�뵚,w��%'6�z�˫4����;��p&����N�~yY&9&}�����t�I�`9�����X���S�!�NE��z�ʾc� �C(��9&�/l1X6q�%�Ey�	��l���S�w9���*�֕�U��2K��`�*Sn��O��
�7�rػ��.|o��|+�rh�Xą7:/���
j>e��8ڛ�{��u/�m��a[�3��y �����A4TK'�r3EOK�o~b��t���>��p�2�����'�Ja�L�樯V������H����,���d
g*���e�D.�*�����n��N�(<��G�(�����@K�ohB�NM����nN[������;_��o ���U�XL�^Rc����*'�6�){���R�֞��9�!I�e�O�8e	!вW�#���	i_s;���)R=�Z	a&)K��xI�YK6ۆ'�rx���6,���0��5�P��O枵�����D�׷�i�4O�yS�I��� '`���i�<�W��K��g���H�Q����BLT�z�b�3�1/R�Ҩa�G��O�9�ҳ�o����n��Z�����P���m#kB��G�lM&�Rhٖ�r�<�AI6�ʟO��&?
1֎(�w�Ecu�V��-��DL�>�)�.��E��9�]�9:��!��Ætf��G�[)n\�}�GN�_��8ڒs� H�xg��:�Y ����j4���2s��h�8��3��i���
L�_FD͞��-�RWV��7�r�A��H�w��dU�H/�zw�8,z�oz�����j���(Y_3i@X>q	,�[��ٺ���2')����d����}N�0��z���z�oJ �ݪ�U�)���0��i:gF��Z.9����ކ�KunۂքR"q,�:6}�{y�i�tsQ��Z�y�ٴKO��K��:��_�,�\I�zs��s}V'b����Am����I[TD���>'	������� W�	����"��䝚do�8�$Xw�(:�#�,�ݢ���3���V�@fi��^q ��T�����X����ݫs<f[sr^^���Ի�؛o���i�..�8�tb��M����=v懲0Qy�O΄�N��)` v�6<�����j�9�x�ݥ~rg���L�?�hm	�9�r�m���\W6>�A'R6DiG~=?۹�'�<�|N�ŸaK�2�3Us	�����,�v���Y3�5h�uG1�S}]�0K��G�o�o.�"[��U�������P�3�>�60�0N�g�z�V=G�)���f����%*r2GLS���ЭY��~z������(����V�;:� ����ڥc�PE���s�:2:��e�#�-��������%�;��E���޶!�۵�Ʋ�z#YY��j�{L�&��KwxJ�/`�l&I؎�D���S/��tW<�����w&�Iz�l6)t�Iw���dRE#V}����:N��M9P=��S)΂[����������"�[�[�- 	�5�����ϰ�/i��]%�N�*�$��j@�;��c��:�Z�yB�v�Z�\=;��㍽����O�6෩B�0��4��A�\߿��ߺ���6 S�a�(���=F��t����g��3Ih,�v�:��R=L!��?X"��C�0/U0[��Y "N��݂�l�XU.��0��j�O64w��~�Vk�����Dy�aDt�jD�M�0���R���C}c�����<��}l.nY^���J@6��e�P��G=a�K�k�ݙ32�H�Sv�@L��Jr �)���UH�qv1��h'c1쨠�]�2Z���!���z�f.{T�6��2�ٹdt��B��భ���θ{�"0R�=��i>2R�ܫ�m����?�f���r�ҽ"n	@��9<�0J��4,�
M"f��:���+�M��2�0�;w�����N8�x�V�T" [�l �
�r0�t �%5ܲ��N��1��>{
�����x�)��u�2�w�������] W��4:� Jvc�I	H��D�+@������9����i����|�	 5n���i|E�4��f3�pp�	���^��P9�d��*����r�L#;�����tI"����P`-�+��#{�>IV҆��-fuoV�\�N%
��X����V&!y�y�"�Kx_��%@���=��Q�<�{�^^aM����J�=��&M�f���v�-zh vC�� )�~8A��(F#�էI�ˌ����x�����}�v��Ws���`�ŬJ�W2?
,(�ˤ�OA��Cr�u���ޥ!R��h�aR��b��o�9sJ������G�E�!�u� �_xS����F<=�~�I}��>3.u�Ju�f��_���n��Nc��	�Dt)��������� �Dh��}c"�	4���ʽ@�u	��7�������4R}�@hZ"{�!�9�&_,o���v�z���D�Y�%����`U� 3��cK:_C��s��L�X��H!v�/��)�լ�]7q1W�^~#�𭍲�������`~����v��s=*�1!��^v�T+���n���9�q�:�bqlzt�,�iw3�57�� +ॲ�C~vmyI�k�F�s �������:k�u,Ϻ6~�t�E!.If0�J1?k�"��]$U����#��t���"zR����t��4ܜڬ��1�mD"�w!�����`���𒮵��j�@׾j�N��� n!�Ư*;�%�N���aq��ώ#��ڶ�1���\�}- WȾ'�D��̠V�a̺� ������FF˺J)�R��p|K�P�`x�9��
0�XS�9hQ�[���<]p�@���B%J��k3��H��SK/K�䷧��I��Bʺ�ήCu �j��P�Pt��l½K����c��+�ZC��Y���44 ��<��D6�Jl"���|^D�Ү-$o;����/V��6�S�~7<`w+�-U8j�%n��2�C��o�u!<
G���9�d���Tg���om%B,�����@8��SlW0�2L��I�v3�v*�X����κ�&9뀠o/���G�����ܦ�� �	���;�}ۊ�x�n�)G�cl����� ~\k�t�K�4�j��L�`#=��Ye;00�|F�N�

�@}B�mu���i�v���@���tکS�����\3�-�QGA�v��!���%?���>�\�F%Mёo������� �;�M��5�q!+��<�E�	aE@����螦c��r�B@�ϻ��g�2��tL#�O�W�&���I}D��?��f"[��� 1JC s��%�d�����T����i�ʟ��!|X�޸]��r(�Y�>�_9�A>���+����3;jo��b-�Yf�\��!�w{bo{���ߥQ��x��7��4q���*}Gb�sC�+ѱ4��"�8�k�DG������S�/Ҫt
e���.yq2t��&P�[}'^�|�n4ݭ�J��ޭ�6t��O���_D����nX�R��h}�Z��+��y�Yv�У�z5���3�p���h��)!
1�[�(�us���R�EG��"X���z��=I�Kx�$��ý�g9�V��T
N%�����h�L�w��_�7�Dt��!
&�����/vT��چ��q;]��qZ�\[�!��M��FٔO`�o��U9�l�f��oI��O9�].���;zL�a�WM�={�x�Mb��a��B�j�>��@G�Lk����(�M3-��"oV���n�)} ���Oc�R�+� ���b���3�ȡ�80��H�1&$���p#��HM����qZ"�Y�g�e�bB���Q�Ӷ}_��UH{�ս�"K	���D� �;7������sE(�Ʌ�핂g�n��;�W�ݛ�wk�Y�iD�d�L��r�J��q<��Ƴ�$�J�X8k�M9���?�t�J���cB'0�z�\,��
��o7�ro\�|
����b&(J��>��2�<�T�����	�u�JyߕjR�z�u�b��$D����3�����H�n�ǩJ��D�Xl�&�w��1�C�<_�i��?����o����b�J�43|ō�<a��ȴ0��gA����X&��D�#�5�*B`[d��y�,�a?8�J�����B�R�����g�'��s5].=�K�o,��u�ӵq:���V����&�:g�A��TT�G"��?�^ޖ* S��zHh��w�1�2ޙ�tJK<L����s߄��� �b1��E���'.>e�����Ó������63CR��)��+�nt��)�Ŷy�2�zrjX~x��������G49j��\�=&�աK^$�HpDh�����=��5u�����9J��Y$���g1���T�M���V{��Ů���	�OKs��ג��|��Uʫĺm����@�Afu@�[*��`�?UF�=�D|ڃ�gؽn��a#w��dl�Q�i�P^���ք�_�Y)��qU�0���tDl��y�YA�QN%lvSG��l��P�`j9*w����G^ ^��A��g��Ǝu�N����:�z�^��E�W�$����PA }ă-5Drai#[b�{P؅��FP#<_�$35~@�_���M6�·�$�����#�먀@(Iu|�m:����=F�ÂgJ��7|QR0΍j>F��^�\�˒X�,2)83B��o�����l��;Q��F0��g�=_ o�� �I� l��v�t���iKTE��_�(�R��1���"|���, �d�Ad��{�:�G�O��Kb�����.����DrA�OjoX�`p��2�ɶ��-r�S��#�A�`���ޅ�a�������#�9Aç�D��
-��,t�E�L�bz�j9w0��dFQ~�	����W�
�DMO�`��Х����ϛ�n39���X�(������-ą�qo�w�d�U]��K�	���d�va���R�4�HCs�Ǉ[���4�gwߗ��Аd�ݖV�%�F:�Bɣ���M/$�~�`��|B�@�sB�W��N��/�J
��w��*x����ps�b�p,nD����-2��0#6���ޛ��������ܪ������r7G�o�,��_@-9�e�}ֿ�baB�4]4Wb��ڟa�h��p����>S��FX�_�B �(6H���K�Hr����f���r�U�:ku��[�v2��'���i��؂-��ӭ�g<(m��y��:��g8�6��%=�z�¢�jĆĜ�� z���ŸV�@�>�"����_���L6�W��9����U��h	?HW����;(�(���Xz:���[���\4��.���`���a=�a7	�u�r�A��]�aʠV)�o��4@ ��_w�����F<4�ā���0鬃��co���B�,�����n��F�Ad���˯�0�y�\�y�@"�����jnpY��1��E�-$������z�r�S��q�ڢ}(��[ڠy�"ޣp���{�w��a]_��qʧ�h����Hv;-c@aQ�Ϯ�*c�#��z�������xsH��MT;"m��"�t�J��I�tA�~d�-ZU���~2f�p��xP���S?�1��q4ZP��a���oU���C/d���j��3�~	Sۤ�yM���z0�_A��wB�+G�j^6���������f�������n^8n�`�ȮY0ͨl�*N�C}9���/\|&�Q� ���ό`+<�����t�q�\�x�n��4�w�q.��?�]+�6 �,���G��v��� �ъM����q��ʍ���lI6�������L�!�Q7�zޒ�ދ�"T�D]��c�|��h1ja쏡�[	p&�b*=�	�;��IX�y��e�5?�!�'��awJW�{�&$�'�$c�dvu��S���w�u���o����d�:��������\d@S/]����1Įssj�ĮK���.���e�|CG��Sb�V�r��� O�11�5H���t�����9ω棸_��$2x��ǓF3�m��Y�U��2rHA:���}�D���Zz�L1�XK\?9o����4���KĔ�����SG�RYG��՚-��������l���g���C1��,���;lE-�]7�r)�y�������Q�h��qY����A�Y�j3�rŌ)��x��O
���h�X�{b���[l�G47M�`>�h�u��R�|�L�#����O#��⶘�1n7	�����`���\�+��>_�mf-A ���v��  qr��A�:��ց��,k�D�~L�c���!3�����geߜ�f ��տ~������D!kY�i�����pn�;�;��6����h��`T�j�T3L)8�@b�4co�s+�nIf�F�Q�f7�xp���6oLԱ&Vl�#�����?
��{6l�[ �s������sg,&��?3�	��^z\h��^F�5���Q?�i"�w����]68g�|`���0%���D=�rk TF��F'G��>סhR1���ip&��8ڙO�����!ڂ[kC�omA+����Ϗ��,�K��l�g�.�ְQ���r~N>���O
�\��պ`-�}�Vn���g�L���<�g	��b]]ΗԐ
�qe�F.3�S��Q�)S�3h�_�s��5>���7"�K��:C����VW@�á����c���V5�J0v��E�JCZ�A��V�M���4���������_��.	P�Vt~�{m[l��6.���� ���l�R�ۼ��*�&X ^H6�ա�F���ځ���˹����#W��^n�s�ىR�:�+']����q��!t%)݀�;	�'0}&sRӁ��"v�򸫇F[Ly1S}���:��f�U=����MZy`�2�Z4<�$�����G9۰嶁K��S;�a2-P���{_I�K�q:�-�]`o�������(�P,����ˠ_��ի����_i���}̄չ�=0�ϖMg���� ��ͷVI~��=�.��eE�i�����]���#X�..�M�Z�W��\�N�u'DA>����nx�A���Y����B�|��i[|x�Rb��:�Gj���z�[��2|O��&_ȇ�Q-��̢tHG�]=!+ ry���g&���������$SUuCI�����O�>� �KJ�
9�r��I�L��o�c��Rh�#.��g|����p˘+����$��3��-�I��@������(����6"�я1[!L�8nY���5۩O��ؠ0/uc��e$$��衶.��8����Q��ZV%��w�a�Ƈ��2T�	��N�by���dtH��!]��Cڗ^��0�3EF�I�$c	�6n{/�m�3M����Fen�^�^�ͫ��a��r��y��.v=��KE���f��$&�(H�,�w�P^��.��e�� �hS���KF^y�� ��e����H���ٴ�s�����^��w�K,�|��n
�oE��XR��w���_:'�2u��D��� Bx�|��N-\<��z��F�j�ćO���%�����ٵ��*���a�/3JR�Y�}cJ�xFU)�fp�I)2���>�<��Hi�'�����R
�{�Tƾ��x�nlX0&�$N��x��ǵ�~��n��f(��XX���t����k�\T�p��\��F�aY|1f5Ƌ������_=L��M�F���;��<֑�mst�U�"�#��m�/��f�-)��ɠiG;‧�)�K�+ ;T�u�#0gNk[��O�z	9c;��oX��&�E��_��f�4�:�����Y��2��d�\�p$ҁQ�fl�r�*��#/cj�;����%p�(.;R*�1�A���{a5��x7�4�O�]Ȋ���"�./��mvJ.����InCT,b��
�X�C��!���a!�:�ǧ!f�C;H�j��[�����^�ļ\���hj�!l1���Cw8x-�m��c��v�EAe%��S�Q���I+����TĂ��+%�� �~����6D�:�՗�ݩ�ŗ�:L��l��q�=�LK�|��fA��Z.=���o'O�;G:�|��v��Wp�����HKQe�V�êq���~�s��U0#|�!�c����dB��2�~�2Ž�����V�O^�Gf�v�?�g����J��EUv�{��nw�
<�z�@�!P�D<��ޗ���y,h�u�$���+p]�y<	�����m�@m����^]Q[���hLEa�`�v���\m�
@Us9b�6LOW�W�2Lh�I��gꭠWB��S<�=��-�d���	I#8N��Q7�A��8�O9		x~�[�\��):k[��q�x�Z*�����`>Q}T��������.^�,�n%����ˡ���]�?��*H�Q�c<�����}LX�&MqI̬��j��_P�h��#��c���aP������O7��I��\��岝���|����H�������)2$&�z!J�3�	�༢טX��tn}�4&�"�vO�@ہgm�"?b��TqR��g���+u��U��{wm(3-l�&My�?*Jb�Y��R���Rg�h�)
����|a�R�PDxb�	h��jr�?�X���-��Ɣ��3u���n�F�V�h41���#ǟ}tM����ᐎ�V@�Ͻn��aH,�(\�C��(�Jgb4�-���&����q�߹SQ}[;>���n5� _c��Ωz�m��#OE��ÞQt��oU"lȭ��c�A��D�e�cyj�-;Y��SQиm@�n�Y8�0�����đ�X�+LT����q�� ���Tק�ܸO�ỡtP3N�BT�C`�%,Š! 6�/ ��z��ǟ#~\��^���9��;��C<��@�m��=�\(�-��γԥ{�E�4�XN�	OHݝ�f�Q���x�W��)���hǐ� �Y�4� t��>���d�TP���(�j�scf��uW�|I�$F�\eK�Dr:������x�	= y�ICg�ƥU��}H���8H�@����ć,�~d&��`J�U�� �_�1��)�����w�9��5��7�M����d2��A"�k�0��|�h��T���M�_�'��H�yD�2�c$˶��`�h=Un����Gm� ��]P�	ݵy�� N�U&��nN��V�~�#�n� J��Q�&���%�3�2��e��'�l���Q�UI�>` @�l,��oZ&���h����+~�#� l|�E�ܙF��B6��x���*P�5k��T��0�S��"�9�ؘ��e"<%a���x����_�/M�v���ؚ���2����q��~�4��az��u�纊T�y_W�&�Pꫢ��/}:�~'䢶��#h��yOt�veȈi�91?��<�盳���?�l�,d�F �*|��%t���n.jv���P��N�/Q���CC�d�B�c'��x��?O�v����]Ĝ{	ִ;��@8�x�s�F��	��B�qI�6���5IF���՗�n��X'��Q]�|�DH��y9î�6+_w�a�Z�N�4���<ťh_��Q�Q���oM��z���*X>9t��P��r�,�� i���gE�uxw;M=Q4?U�"�����ҤVU�ЉUm^��*~�w�����U�ȗ�ؒ�	z���$�m5���<�,F��O�zc?�4��(��?�d����&�GGi����/��.�)�L=7;�.P��X�v��m�SI���w	��N����9!w7y�!�2�8v������7���o�jC�������G��s�V`m�����kjч��2�0�tj[�ɨ�!��Bp"��B��=Xsk��A���7ɧ<(����;y�^ ����x�J�O8�i��Z�T����sF��Xg���'+���c`����D���G���0&p��>�8_?���x��پ��|K�GQK��6E��z���m��md�p�K�E� -�s�'==����҃���mY�xTcB2���>ב���B[	���}{�B⯘2����Xf��T	��~I^	r��a��ـ8Q0`G��׃Ӏ|mOU#;j�y���#��k���q�R>�y%T*����7٥��!������ ��v�z_�P��6#N�W��Z�<�����D�̤��P�o$��1�Qqc�um�ra4M*�8�S��4W_��i����>������v����
?b�IC���mR!6ie��e���[�Ɇ��ٟ��|:@܆Mܧ�u^D;k��q���/e���"��Q��b�P5�x��(�-�ܯ� ��/k�:�Y�)$����فιG�ڏ��ru�!s�/Ƴ�����۬X�ׁ̈́ a�X���U�*H�%=�>^k}]l��=�J��6rI�D.B� K=���+��r:>�'OH��FU"�t�I�����1��W�e7�o�%In\9ֲxA�Q�J��#�%�|�:ؕ1>>���w�#�#�|���Q��������YU�p"j�|��1�h�}ـ-��'�w�(�O��Z�t@Hl���RQ��B	;�fA��?+><�{�蒠D�qh�*�w"����u�M��W?uȧ��+����K�c�͛�Y=�˟-�h��LV�f�=�+�H���#�刌0}Q'#[�#�&OԷ�=h�O��<=��Yg�������`FCI��2/H� ����O⺦n�9�����G�bL��A�����چ�,G�_e�Ѕ�8F0j��ˎ��`�0�M�`&i�GMm�;.�����C���q'_,��=��=�j�P��G�B��)^�\	�\��sP�����{"�Jgc��WA��!�����*��l����`���
"z��u�C��Y�{��VYA��v��d��S�ઌ3���d���*n�$��U~[_���O�����/hGG�sb�N$d&�u�6�Vţ1� {�V���������"�
�,��:�l?��u�O�����arS-�r ����	��_F��Oh���x�}��~.;[�b|*�Q�x�mry�Y�!_x?-<��9f�*�ǅ�񙅅(3���4Q�1?eIm�R�#Z��o��d�����oB��YͺJ�v��v��+�DI�d$;�^�\AǑ�UĐ�����0���4]V��7�9\r�n���9�XK��t�1���c���F��[Қ�Y?�8�a��0."�Dɛ[�9���Z��گi�}sS�SA�	L��&�o]�L<��J�Q�ǧ�� �0v���#�<k�xk���A���j��u.R :S�b`LNH�DC"�	�*�14V�噭 A4:T֓2T�5�sC��A\mKaϺ��Y��Ч� sJwx�a��Ig-�,�!S>���4��^ys�|�]~e'���J������_�r�=hM�pu���;�����[ܱ���d�ṅP�8�dF�Dy��JS�Lc~�ȕGO:��uE(-��/Ꮤ�7_��6�w�no�����U�$��V����83�x��l��Lv��K�����ǜ7[���� ��O�=cn���#�^DD��<А�-Ti���%��Y�� �<+�m;	QȢ��L~�"_})~vH�~�W�,<�ⵑ��_��U��+�R��b��|CߍL��sɣ4g��{��lpkMC���#��G��6½+�J�T�
�V��w����/`;F��v����6Ks?Y�8v��[o9IO��٣�V���L4�Ñڥ;�X�N�>^~Rx�ܾY�5P}1���}xT�1̆��ى�P��ly4<G6��`N�@	5C}?�>�k�O������s�T�8�Dꯦ�B36�$qP�����7�=�v��bc����(�k7O1�vzq�wH��U�D�Pva��� aI!��+�.O�ņ��X+�k�a��P�w����t���rwi��h}����G��4i4P�F]iw�u%�%�0\�哥�e�}t3vA� �L���d�(9T�s幬��qh�_|/����P�����Xܓ���܍�*Ps)_D/x�����I�S�
�z�2`��7͸�+���˓֥��~+�}U��#72������<`�v����n��!�l���HD�M������x�o	��*�B[}����:[��'�6%���h�Q��F��G�����r ��ۋn�f�r}W�fܱ�e�8�چ� ���a�1�,���f*��mR�4(�i@X���7���#x�-�\�d�A�X~�i�]���Ĭ�cjh)GynB��n�&���N�I�Ð;k;{7"���?;&ރky�4���;-uJ�����?h�X�4o��W?�eB=���^e\�;{_�B	�%��9���m՘�sd3J���*�w���Q�J%�Ġ-Z�q��԰�̝�$���d6��[X�;�<�.��9��ܔ��'��7���� ��l�>�~=�����Q�@�Z#i1�@�TuK٨�C���+��OB�U�����
�����gH��t�.z���<����Y����{yKT
'�3>K4�]޻,W��C��'L!p���	�oX�6��$!���~�։���(dGQʣU�.=3@|
6{*4(+�9CDSV?��єȓH�����M�S�k<Zj��∞?��>ahx�|��j��=�f�e�H־lN����ZL�`��s��v�c)�m�;�����p�eG�T�o��)����±��K˴.����-3��4c!��@ ��|��]6�a���^}DS|L9��7sqM	8��VB�+ TO
U��ټ
�Sh שG8:��jzg�g#l4�G 5��SB7�>�s�j�7��򜴽�l05����0�� ���,�$Ky�ƙ��dx ���d{��r�0I&uS�׆Ԫ��#@A�Dp��e�~'��pC��~5�]T������✐s?�r���_�w��*=��P-���x2�X�:%��k���Z,h���Z~xM�R}��f�O� �%j!�3��DCe�$���r�����T�R��oD:���-������`�*&pz��XFp�@+������o`\�bx�BZ?��AL�C�K����H�@�^��}"]����H���fa�T��*��(.���>@r�����B{�qL)����u���]���9�(Hbi����h���<��#�7`�D�ҏh`��*��K��˨��!����tZx�=Ơ	t8CvP�2H�`�T�
+4��H�Kh>��Lc�hx��Z��ã�;k5�s;{�})���Wb��A)<F=&j�$0m
��w�t�ĺ�x��	�lM���lt��pu0�RC0v���9��yġ�`MiO�l��/�V	^ǖ��uP�qq�
8FVo�`���Sa$b��3�|��\���9����e�DMBAy8���s�o���Y��M��JАf��MiNX7(҃:�6�vj�	;^���G �X��Hv�"��e��{�S3ii�ҿGp��Q���wBΊ��S�,��||pb�/��#N_���$ӳ�bR/x��3"#dwB5h�Bl��+�O���T{��d*Hj;���%��<�M������`d�~�!�������K��K�՘�U[r:�2�Ӝ�6�L��C��KP���B�����"Y�5Ń7e�H$�Y?�C��uH�Exl���Q�_ΰE��~6���o����k�H�E@QC�!�^��hU�66 k�m���#��o�碲�c�/��gb<�Ezy�H ��a����z_\4�)^LIމ��>ߝh�+�1�Xx�R�j�h�ʌ^���W�F�c�ϡ'Ng�?ۻ̵輿�����~J��#�l��*��I?���4MS���o���d;��x�XOl�W�!l�o�����Y>�0?�:��ըAZ{44���/kI�uj˙�N����=WTƇR���ǽ��G<k.��C,_P������,-��-�K�W��y-b�2̾��4 �i�H�L�Zq�F�T<`|�4K��î��2
���t�{��=�8��S�=ND�#�"�C03ݑ:�25�Ρ�1M���@�ڭ��w��f�BI~(A��j��7݊�D�^�.^��F�G������]N��ģ�"B ��chW����~KAj��Ѯg�4uMS�¿2�P�)b���gƻ�E��t�L�?� 3�&�<�gغ\҉���v궜�T+��v�	�A���J�kRzB*����c>a����<\��B�6N |w�Q+)�6��]��(0��%��*݋z�p���R+��)C @�`�o~f;���Ӭ+�z,���*?-WI�"Z���8[�Zq�P'-��9Ơ�_����I9"6
A��j$�C�3;'D�r����{��oc#��z�^,e����V�oU�����
�߾T�]-�x��S�f���Rq5��SH�k�׼Wg��v�h}K5�_�ܠ�y�TK]D�p�
S�k�nW��|�`_*�-��D[o~B.�Ϗ�+E�U�����5��h��*�^��X6�#E#�5(���:�s�	0�������\��!�x)=��^c'k�)ж�֩v��?w��1r��}�6�����%��4�I��6�-�E�X�<����Ut�ׁ"�+��	��UD��hڨf�/db�!���Fw_b}��W���Rn�������R�@�:G w%[��GK�͐f�
�A^g������s�d��5o/5��U��~�Arj<��*���i��f��}�ۑ���"{of���w�pp�/.���p]z(" ����~�6�BD<Բz�9��!��D�5�i!�D�ɻ�I��ȱG�k*��u�|o<�[�CG�&_��s
c�����جY��M'�m���Z! ڈ����i
k�h/^Y�}sc��?��_&��aa��0'�QR�8W7�z�Ҥ����B��[��=/��3���΀$�+>l�_ AhF't|R��OI�t���nգ1S�A�f�_��f���fsǰ �ə���G�NT0�5G�O�O�we?I�pU8���'��>g%���U.1	c�>,����k�'d� r����i�����c���f��c�T<�8/F��b�'\������}�f;���<�)��Ҭ599��s��ɀR	�ZIW^��d�[��,�U��Cg,�0)�"(��HΠ��b���y�I������>��k1�Yܞ��hW�r�?QN�(/i�A¹��g{���	�p���4q���,dD�/�$*�~O�/p6�r�m_���q��2T���0ex����n��,���Tҳ�!��zH��.�O�Axh(/8�FϽ����&
�PzWYD${0�x��k=�d��N��?�I$��g�I-�xM�q�
`�K����3�����%�bh(��mT]aOӎmF�՘�9�ڹ�	ʅ�K;�0��FC�1���u�j ݰK���*b�}�+V(Q�B���~<��~Āh�N��s�ԏ��Y2Qs��5UpN_�,�zWܨ�{�Ao;s���bNM���I!:&�nBBJU-ӑ���Q�Q�5����,��[��1]�vM7c�ƶ�a�La q���L�=2�8"��0h4J��#6�R�����M�	1��J.�D��g[�q�F����h���%���S�a�%�P9~�U+��p�7F�b�.�fW������>�������Hv�C�K�8��<ۺ�ճm�(�Lq$������7h�≂Bt59��x��c�L��,�ҴnFl�B��m�O����9��O�e1M���[д�b�"����K�GS{���Yܯ��
4�0�F���f��o{���Ǔ��5�c]���L3A���e-,�Ih���mK_"��9:,��Y~��y݋��vP0�ߴ�޿�f$��ЦE��y,Z2����e�T�0j���5U�E�s��D�`�kZ[�_+���ˉ4h'pH\��1r�4�űӶG�/��'�?�ӄ��<��������]B�N�R���Ջ*�>��A�#ƍ״:8���i5���t��BCU��%"1���˸����ȖK�'�y?�s��ۡh����!/4���oڔ�"�!�ư����iP�W����3�ĩ'}�;�O}I���:[����,�10�P��~��=���{j����H�1�8ӿ�3����W/l��_���c͝L�g�+Oё<��*���vg�5�����J9|���b{�hxK�V����y�{���������`�s���L|?�*��'T֘R/��@j�+Y�8Dv�R�*ɣ"e���h>��c%c7#�w�n��xVV�o����sL8X6��M�e;_�;���ACBv�:� ��^��W��v�X�?������x#�ڇ�S���6���`�_�%s�N���ox�e �:�0�\J��H��I*�D�P�A�l�]e����e�%�h����bͨ�*��xN�F�ad�9�H6��j0mqj|_��k����m;f��4��T�&�Bʇ��|2�qr�X���[
�h�I�E���p<�>��wq 蛊���8�0�H?�r`��1� ���.��w�<'��u$]ː����:Cwճ7B�y���P�-���ps%�4�f8��l�	!�̘J���g�?��6����si��0���o��j_t�e�����$���� +�6 ���M/f7��ZO���3y�WTFwoX{�Ԗ�t-E���4y�Ѹľ�1, F�A),1��F��4/���x���_��Ý�A.Z\�Ӄ�G����s�=�v���}Q�����=�u��':�Cy5M�v���-x2��B���!%%�o�\�\Ak?��(Q�笌����x;�u+&!�V�����L�E�����y�?�(��^� 
X��'� 1! G7y�XEҭ�`���:J,�B<R��D�0=kO��bC�����=��<�f��3�ZRf�HY!`��%F�|���\�k�5�KO�(C
���z����o��+��m�j����B��(&�O�o�A���Rಬ7�8�U`��
�S��V쏘D���N����bB/��(W;����2J�a]�nQ8�G��L<OQ�����.��>��l������ܐ��@���I��VUͿ�$i���3��F�����#�<����Q�65{6V�X��T[�uG�T�g$�\�)��g�5i1�>�u���tl.�X��昢��1���� ��ƙ%��k�?W���K+�{[�3��z���	���^$�E��6��K�]R2�3����*j�q*�mo����9#�[�� �,y��4��r����K0I�;%j��Do~�nF�nߥL�E {���?d*i� r���Ǆ����Nu�Z7V�q�z�����C3�J8�],�RZ̖۷+�V	�0�L�:��Ixw���LɖBx ���k�k��H'�+3a�R�W1_xQ	d����h�i��|�e����\�G?ǍY��^�2���;��hN�K��7h���`S���s��&�>L��v�$=ʔ�ӃO���=�(@FRE���t�!`ۇ޳EҎ1/�.>y��;��� ��f�᧜E��l�
Vڒ7A��ГJ�^3��pɆ��dM�~ţ�����	�����%�n���q֦����i�y>7ɝ����<"����O)T�-�(e�l`O��<-ݻ�.�_L�������e6V_s�Q�g����x���vzwT��!�K�	.���J�:��$�DZ�uƿ���Ȥ� �`��Z~��<q��灍}�k�6�'Z*k��	'��$=���ˮ�b��F��Ţ�;���G+_�3�s���P�����r?�)�A�J�e4�0��4�ۄ�r�UK�Ԑ������e�3�\;�RJ��{F��ޞ�]�Ѿ.(i{���G� �z�+���B�ɷ�����x���Hu�㧙�Y)�s�-��f�����i��WX-0�$|_����eJ��^�����W�OS�`
e,���aE(N<�Ǹ����T����ص�t?��֬yXrkko�a�V��w�k�iف�gH+t���䝡��~��G΃ZKJ�g�w��gOV���M����i�>�i�-�|��<�}�C���'�թ�`�7H�DcnA��3P+~����e<�.�l=�j$�Wܔ+�0U�H����+?������`"� ��1\��/%������K���n��Of��M��f
�'����)D��m���ŵS-����-��,��֫��k��E��/&��V����G��Hf�=�e��P�մ�^t4��Ľ�����Y?RnQ:�֬3�Lo4���:��nQ�������`Q.��@��=��f����m����`�i���#|Oe�,���U���<��a�������"X�I�Dw��yц���2���;�{^�ϴi��JI�����Oz՝^����9d@���wVɕN��l"�䆯Fݑ��.;��Pq&흯�8|Zxq*�Aߺ���Suۑ�����^��ѯ���g�_/`���(H	��k��4����w¢ mP��y~���4oٟF�F�������Y%�8ɵ�J�A�S�lVe�+鮤w�J�2~#�X���,�^����țӗ��xW��w��9��*�*�,PC�+�=,V���#�L�f��Q	�=k�����̴�Ca��Y�󊬌ژ��A:<X��\�9������K��;�a�W�o����ס��yXF�|��X�!_��J	�yt��=��|���q��W1#�- ��;�2�܄WP�����F��_�]�'V����U�������Zm��ϒ��Ը*Av��_�0n���~Q%ް@|�_�{����ɬg�|6�W��i�j�5}�@f�sQ7
�����W�u���u�"!h��pqK�U��sW^�22R�a{=A��
�s�����$���^���9����-� :A@�@6M`������۲8�Vq|�վc�kl�B��v��,���A��܈��]O��hv����Μ����� ��(���^9�ْ'�&��h�D0�*����Hgl_��ܢ�y�K��l��t	�	H�{y�h~�wCe▵����ߐ� Ћ�}m��틖.��閾��� ��1�8�ގaA��V"eJ���c�m=+z_j�RB����I��)����A��=�����!��?�|~¬������Ïu���1�dj���K���+MK6��u�ູe�l�2�Z�拣f����|{�޶OH�6$f�����	g��wIS���Qql!��8q㐞�ҜMv��b�����7�����T����� �xڌ}����ߦ���$2�C��J���Yړ[����ރ���2�^[	�1�����i�j�����O��4%��/����v�C��+ñ]Lxo=�����Y�y�~�ȋ/�n�"@dU	,p��A$6_���G�c���wv(�h�m������� &��G����H��	 [�j�S� S�ј�i%�ƶ8�Y�O�R��%��x���Cg�R@���2a6�;�
����1���{k	����q���lGu�7V0����'ۋ* ��L��2�$�T�=�Kљ�7U�)��XZz�-���{�t�a#Ϛ�k)���j5"-��-���کrs�O~t;���N�r;d���(�Ħ�G�R.M���Ð��mqN� �,�i!9�`��� bl,M$~͎�&M�7m�on5�G�B�n� h-*��9ɑ|6� D�iJ0]�Ǥ���B��.Uӄ�k:0�=�Pao}��f��(��F)e�k�6�6�r)���`r(F�S~��>P�a�\��E�H�����ʎ���vI�_H{ϥ�#�D�c���w�}��G\���E =?�yd�CWL~du��ld�ǚ���$�W��He���9RBk���F�e�A���f)e�_�_m8�ȰF��:�!fxW�nJ�RJЦԪqa8(tF�q�:#�q9M��n2^㱏Q�q)Ȥ���xϑ���o3�cJ�1Pm�ir6���=!6ϷCX	˱��6W)���M����g>�ǜo��Æ^� �8���
t���`o5���0r6j�-4�5��|�?,R^E6�{{����#���ǡ7��3�����pܴ�&N9��mY<k�Ɯ��ip%.X&߽$�1�`~H�����T��8u�u�U�M��;�ϙ��zR��d^��"ZYǷ�*���Y*�ܞLλ�P��<�]�֤S��KO����y�T��H��;�bh9J/��zk������H�� U d��F��Y=�?�0,?0Z��ݝ�)[4��Awl �� η1���q�#y �sj�5��*M�*�Ӡ���1�0C�+�����>�y�S���d�H^���]c�9!�����`�5-H��^�7uU]�S�7g-�K��2����#Γ�_+�p�A���\M��K���C�㌔9�8�%�*�uM/R@���G}�U2̷�UIR�������6��l��d�i��wio��-Y��t7�����ʎ�)X�KH<�����n�Sl�QD�I,�F/M��\����G�n��?~��+�-m����{~W��+KN��KH���N�K���8�iЋ��$J������j�3��fl��Z���;�Qe[@����|�e/}:ڒ�-M��E��*V�^ݙco�� D�6��P�!~)�� f��O�hC �l�OE3̉Oc��)��?�RD���l-z�`bp �t!rB��k��y�R\�Vw�W����y�
$�lҀ'����qLE�H��[��1��0s�n杜|o��#at���=P~O�n��7�������*}?[%R殯��S��j����>ؼt��I <R��DgJ,�i/�Iw��U�Mi��,�ia�?����:(��t��g��$썱�g���'`��	�Wg�4>�ٙW�t~�)��(Y�3)n�h0#8$����[�^)q��~�Y���C'~�<^�&t�r�5!��GC�c8@�](�u�Z9�˲g�̺�l�,��������K����>�O����c[���`{�fw"J2ox��TP��d�rX-GRq	�&MO����[��Y��2��M �q���*C)M�xK�C���C萢RF��D�ч�]Ћ���H��PW%�@$:����_�aXk d�ho�B�a���_0쫀�[Y1�\,�]�2�3��pTJ����8%�k���k1A,ҽ��F�����m���	�X��f��~1kOXAw�Y}��P����3)WC-��������jCYm^�����9��W�V!�yǦZ<7�;5AWT.�(�ws����lW4𠼡rs���y���Ȇ�D �ð���*���~!�ڤ��F��H�494�:�;�������@#)ډjU6��a���6�ڹ	����m46$�J#�|�?�1�L�6�[�e�������?����W���5%�?yq��'�t���g�����սY��!�&B:g����%�q��EHqVU��C�b�r~R�|<�� �m������m���Fȗo�J�y����x�:2ҩh��[�%g�g���{SA�{��.�ܮ`��S!T��Bv�b����&*Q�$;��/3g�Hf,������\�}q)�e3��7/�k<����m�"�������4OZKb��������'O�W��Qd���
�3�v�D��be!A����0N����]�?L+�G��j)&�wRQ�bϢ�7\o'�Qh�e���q�%WV9����A�L���\?X�L��h���?dY&&NZ,k�462O�` ��<��z���m,!���a��X��&�7��"d�+���@O��Q�[�.�1�J9Q�1US��[�툽`��'���5�pLǩ�-�7��d�D�u�Y_[�oÓ��;��������nL�ؘ3�p�|�2�?����4`�j��x�x�����RC��V	rл����11�:�����6��OJ	Po��5����;�A|z�t�]�=�^x�N&Z�w/������u��	rp�k�ݫ�+
v��G5I�G#��M� ��w��rvA��ȸ�ͦ�>�Ȳ�w��}>�QQ���YT���e���k�I�v���:);����2oJ�uˠl��-�����ڈ�!��\��rx������0�<�x8�o�K(W��܃F��R	G�M�r#���b9_S��:���ҧ����)����N$����F6������]�� Q~7�>�x\�qY�vʾ&�ś��&2�ט牥�Rz���+f|p��a�k�R�㔞P�$-����0�F�a���<9x�l������ d�~Z/j��,Ť.h��9�{�$�Jp'&I��E;�Q����f��rL19��R !�0Y����������:��J-��k���]M8�oLݻ�g��aöʬݧ�	yj8���؇\�G��?�`�9a�-�2�C�|ض��	n��=���	^���"/��f���r��f9���'6�ϋg�˜���T��ݞn86��c	��Ew75\9y�Е R"�w�5_aMO '�Ewz1��@�_�A�U~��epI!u������Mȇ�L��븽	�2�k�q�fZQ�)\�n���N��n9;$�IQ<䲫�ɭҪ�s��T�b4@��h8e��@
�M/"$9�W�M�1�'IG�vҰm���W����<gS�����4���zQ�`������ \F�ӽ�fU��U�
�6�D�#A�~�\�ׂ}���F�e�qE����^h'�*l���+�?�]�(]YIf����@C� �9gAW)���G����U`�Y�S��ci�I=q�c� ��հ]@��g`.`m�Y �� � R₋>C���(� d�hpr66�C,Ÿ��:<���ʱ.��lFP|���`����.�h��x{8]�Zߊ%�t8J��J,�L�����&���2ϊ_�1k>ٓXF-Q7@EL�Ir��!�����%�/���m�h9�|�<�ή��:��.���swP�ψ%;�
Dq�VZ;z#�v^4��`)����$^0��@�l���y&�Y_A�Yq{��;bK��S=�*�^ZX��Ӑ��_�=Hg�sfm
�D�7�J���i��-Mtl	��165-�n/{�EX��4{I196M�E�c=�@�e�����4V�eGf��J/!�៥��1%����iq ���[�v�Ja�~�dЕ���}���(�Nc���656B��"��^E����ᄊ�~iP��%IOM�7ßl���mˣ�H8�ݎ�ތ��\�B���<h�w�L(!�Ti<ˌX���EcQ��N	�:�˿��5�̹���(ݔ�*��0���դ>#�WR����RV	�����
y����~�3ȑ�d&[|�߅̨�4�L=�3�Ī6 ݐ��*;��.T��259Dʆ:V�zl�@�}E��+����t��Nb�cڴ�y�/��[��H��N���3Lw42�Ԛ���� 9n*bG���0hx�,���M��-y�0���-� ���	�(��e�S}iJ17�Y�G<���Y�0Tf�hv�y��x���Ei$�b�%�x�_�v�-V*d<�"b澝#;����(��x��e2�b��Q���&�~r���2`�Tf�f��[����G�^���}�-'x 2[^6�Kc��yG�����R�?`�Q��n}D���y��2-A�ֆ:�.?��#�U�NyÂ�B�B@�_������f\| OK
�iJ�.�<����ا�~]�H�������8{�����Vv�3׹��VV"�C��Ѿȿ歐"��j�>���H�Fq\���� ���B����z���w,�}���n˗�ћ
G-���q���e�G�ԝ�+[f��� ���T(r�~G9$�Ǳwwp�c)aR��w�4�mh�}*y6�R�X�i��¸������GCr�~�i4� >�'ŏq���W0!������U��º��<(lN�_`6?, M&�AN~��Y�'�J��\���3�G{~���%~�`��� %�}�╢k�GR���\t�c?�����)o�`������j��M�d�DQ`6��Pn�v�q�	9ƀ����l�y�Iη�m�����a��ґ��ID���t2������&;���m�4/I.~�3��s�On�_�a����u�t��V
�R��%y��>Pxxtx�c��?O��@5�Myz�M�/7"ƕs]_'ڈ�c�gѧ݅�5s� ������}��7�9w� �����MӒT��Do�v���ڃo���m[��2c}�f�^�"%�Mz��a�o��\]E���~���w�Y�*ܻ����V�R�7Ʒ����ڭ�}��c�Qg�c4+�3��#MZ?߂�~��%b &I��p鴧��^K\�5�_^]	�]��s2/P����!r죱і������#7���8��p/qR�z|�+��= �C�q�=������i��";����*�� -�Dj�O�#�Q�2l��8�4��I�"����Y�y��pV7��Qt�	�:h�fL�JJ�Y^�n{���
�ؑC*��) "��¼���U�E�hWn�̫#l���.7Q�@�N��cY�8���f����5�g�R�o��ŞE�=�("G�R����"�i�p��1&�dWڙ��5��J�]s���,o���.�e�`�%U:�>s([�f��3�~��:�_DY]]=clxr±^�T� ������Z��O�F�лc��pP	2yi�@y�m��K��D�H�ת6B2hP�^،Φ�^8K��`��&Ͳ�h[¯��@�]AuV���Ɠ6"�Dt/�1����Q�)�g�%ܪW�B���h�A��U����˗&H��*��c7��Q�ʃ��N�_�ԺM��(��E1_��/E:"},ta9Y݅`���xss�)��8��
����Nu	Т�����^�0���"���WN`�g�a�����A�����>��}���s xv,Yi}PdF�^p���]�ˇapG�G.����p^{�Y�^=-��i/Q�c�z+f��b���i�L"��M�TNz3��%��l���@�ݳ�ٔ�,����y��t���~�{1b{KQ�ˈ�徖�z?�͸��6�n��qe�zش��?pg�V(�!N���RU�F�(��/Z�����JIi���^r9�AFY��׾��g��gV�n���PNB �	LVx����ꏶ20Ӆ+��iGC����_����H&+���*^:\�3\�Ҷ���FI��P"AD��Yb\ؔZN�a�Z�m/��_�q�~Y/w�g`��N�p���t]��ҪnM�f�9��%/E#��Һs?�Յ!*�X�kJ�Ү\}!]�G�2�0w�;��p�6b^�ߵ��g6��е��� .��Gf3n ء*����/��Xqs���m��%�T�H���
i���Oї��VV�"~�e��	����#�:+C<IH���S��v"]���	�mav��$rrq��U$M�ڑ�{���E	�s�9��xޅ��~��K�tiV�vS* �:60��t�b�T��9a�7Զ�)�1�����9�l�Ѯ�I���c���Xս��������)MϷ��`��7}����4C�x�V`��}l������M�!�� pG��L�w�=�>	X"�uΑ�o�+|�gW����sބ	7��g
�P���Pff�$&��~�q���<�6S������.�����C�w�!
�޾���1-־ک�~���-�"�����Y�]O����Y~/�mK�����ǘ����A<���L��8�g8<�T���S}�:�xK����2Ƹ�q�}:�񪙀-�&JE{������ў1�0e�Â_�:ͩ�n#VW�1 �1w��2�I5T�嫷�h�ӳE��Ff 7�ENSg��������(���EE���ƭ7�t�h��#?��~���!l|��fU� �j�����v���gX�g':�o��3j1�d�\O׎��3����?�'��]e��/ƈ ����\���o����{f)]�k��p�~����g"��2�kd���ծ߰�^��vx���5��iǈ���U[+R�^��@�T�d��9gu�Z@l6z9L ���k��־*��p�5!�<S��׳
qᏚ߱0W��f8���Վ��Q�1��׃�c�{���e!��c�	g��� N��:�	� ��c3 ��m]�4���Q��h'��O��3��Y��H�z��֌0=��X6`H��(7�A�i\p�d.w-�����h�s��%��8=���|/P�FD�0q�#1p���n������K� ��#�	���Eŏ�P�o��o)�GM `�=#{�ba����С��N5>� �!-�U��85��D�����r��M�m�3$x�+�,����})�V�E1�G0��z%#$d#)J96�Z��R���%Q�V��E�ԞF���Z7M
��IQ"�5+y&���|��/�^��c��>�fH�d�X��`ZH�mx���	�e�j���?�m8
9��y1��S�ma;��ӹS+o �M��~s<\�x6�[_���ΐ%�Sk������X���u:�zb��jip�*Ŭ�}��j�PD)� �AfѶ�+�+�������F<ߒ����8��pX�-� ��Eh���E�n�8\���g��ݔ�t��g9��(���=隀�H��#2�r�r��f7����/� �S�� �^��Z��q_��'#�լ�׹��QĬ��ʽ����^��������(;����|s�1���/Q� ]3�m~7�ē��EL*Sq����N�&)�O���˾,뇸t,�gBhCr]�qrY��s�ɌK�j��ƳR�N�g�'KPp/UQ�ړ�4���sɛR#���X��Ț��˒�$�M��eE�/���E��G|E�$`�ͩ�hg�?�r�A@#v��s?4jΆB�[]��U3h�(��i���|r+R{�e��+���K���d%��G*��\��´Bb�*ʻR&9�mb�� �D�FwHQ��;3P,��[�!�^��V֒�ܩ���������̩��!�_͊V4�4��S���ܒ$2��2�Ū���=�
�{w�d���oP=�������� ?C�Ōܘ���"`���bn��������Oڄ�Ty�=U%l�o�ьX���m�o������*����N��=�`�|�wY�=��-�^��m��6#�|h�[?7���o�����r*4Kį#<�_�(t�G�t��{tCG��B!`��1:���e�Ҷ�lJ��5���o�4��>�$%�B���;C�����W�ɍ��`�nDH�~��Ƕ!ܻ3A�AX�Y����3	�B�DNg�~��R�E�Q\#N����j'fOl��͔;�� �4��ږ>W�f�ÎhKG,��dX�v5A�?�)	�{P��T�"�5P�`�eR��U[�p|�	��=�uO2���nż<
w�{n�~�����&-q�$�Y��]��}sACy�h?B{��	$�r�ϗ1��$�Yģ��zg�q��p~eYl�3��G;����������i��ڈ�<ފ� v�>��"S>�x#g�c��k�dm�EC3�
�1p/�H�!�oA7�VyP���Z�6�?d�v�) x�F�e�D�,I�Q���k� ���C).^�����3<?�3��bI���+���zbH��~!%��(��6�����=Gߠ:�4$wP�/�W۠"p�����ud��wA��n�^�M��Yɦm�4��ԅf��[�aYٚ�#��A�G��
�����!%t���Q^پ�7E��ɶlu_p�[���y�[���pF_�&MG*>��4�3�+Q����Ys��Vr����k�(}'5O.gV�~�'��'L����u�qr|�Y�7ۯ�X$ߞ�<�_���/A��ߤ+tpX3�`�b�p{�u�X� ��eW�0�ɚ,�A��B�I��^+R��2��l�X��Ȍ]%�+�{v���z�<�C,A�[w��1�|��w��L6�\W��Kk���Yy��Ծ�o@z�~����7�p2ğ���/D����LN��ؚI�at8��o�0}em̔w��Z��WK����~�>�����v@�$ش�Ҕ�~�J�ʥr��dH��jҭ��%Z��]�Zy^��b}�'x}����X�@��#�6��?c�����3A�m��B��f��v����l#������=^[��� ���P�R+E(7\o�R����1��t�xBl�;�:��[�+�MH,ʖ���`��ܼ��X7�:=�-����{�5��h�Y��0P0���1�l*�������G9&���?����0z���C�a��E�m��J+l1A7��,r�{֗�YKZ
fc-N`�f"d{����3!-D"T�O�'A�ܽl_B���9�(("�������;Uc�
ߚG����4��GGRM���2�K���Q
��9X}_���_��-�㧳��R�w��9"�6CM��W�"v���:�,Hb����r�4kKz�+X�DO���I�+� �Z��N��^D�U���Rʴ̃g�:�YO���:=ԁ��0�*bKTC�j� �)"��nw�gE��L=^��t�E���S�����:�>ӵ�r�iз��% �Mˣ����m�8���_�J��u�3��D#��I��9Tt��R਽H���<���l �{�E"D����i��K�<��Zl�dZ�+��8�3�LK8�)��ɷ,,|�}TVWP�`���c��+�K���)/��sS��-��2�k\8��j6�d~�\���z�j��7��|�TnD�z��jqA��W/�GqMǍ|z�/V�ww�p'QFf%s�S��]�];��`8�5�#	������A ���5@B��
����Zp��Ϛ1G��nS�KTd����J��6@I-`�7qʙ2�m�*ƈV�=��g/((�x�pn��pYx'�>�%o��hƽ|3w���.k�`z4���Z03-�Y��ad�yDh����ga��N����wrfC����8ſ�n�U8�?�, ��4,���;�H��v���xv>�λ�ؗ:�a\�s/�z�A!�@Z�a��X��袤���Ζp�Mx�\k�l;!��h�뱁���'^���{��(O��n��չ&HH+�B|����eU�f���2�`��`H�։5Jt|�AHu<���%���,V�����������_�D�A^����U��Š���h��an�[#Q["�l���[]Q�9�>� �:8�����ޘ�b����g���t�&:�⭘I+F���? �'�!+9��)j�l�<rK��X<�O��L�����,��A0BK8�f���^qp�� 5���}�@&�y��ޣw?��i,��{R���i��U'����5��ΑPlT��+��N6��{��Z(�i�E�-�`j�·�ٗ��Y[y�	v�W^C������I�kQ=y�>0p�z��̔8J�<`?)�c%���8��71��Z ��D?���c&��}a��U�M��i
�u��\�?uã��#�41"T�rWv�w"��˜;�q�R=ʜ�̖�ބ��_e��Չ>��⠥�M���sf�g�Q����+�[�tq���TȨ|�^�$b�?��Bc�:R��q\���q����Imu�	�f��*0�@Pe��M�Q-�����R1 �@���?�ǻ�o���sx�=�VD-)3-g�o���!�m%�u�"�@������J���0�x֦5�qYzw��x�3_�!��q�#���է����C�ثu�xU��G��Qm��N�*O�Q���^��P	d@P:M���[�"M�b��|��[���I&؜*d�|aݓ?�l���RP]�D%�x�ø	ퟩ--�!��U��Y�;3F��g�cNR�FÎ��+��|�Z�L {&ig�uT]��h6I����S�7�a�Ւ�~�=*���u�B-e������o�c]hG�l*0fE<}(��1���(>������ ���6������3�Gń�=�_���g;�#x���B�6��bъ@�AM R��Bq5Em�Z=�DD�Ey	�8:�g��&qv�^�v]:_��L?���@]2G�	���?����������]�|�I,Z�*�E���9Q�NB����`&6^ʻ-�Қ��L׿���a����CYJ;GPA5V��Z�̚^2���"�"�9�� ! /W�h0&z�d���f�>a/.K2?3	j�ٺf\iiz��nE
��9s��[Ҿ�:^��\�1�9��4�R�qE�i��� G�[F��[��0���M�t���÷j����������1 ��xd4���v�=���$PDV�o�l����"���N]㌈�p?���e���x�1�%3�0L0�&UU����`f]?�&@��存����S��Ү��pJ�I�/n#����P�Ѕ��j�쟡�I�t�"�aL�Zɧ��F�/�!y�W�ީ��S�F��)��O�Vuw�_�5���3^�|.�Q�؅WS(��b�ъ��RHLh�r�WĐ�yq���X?����:�����G����x.GCV�/w�t�1�qG���R\��X�\������@�ߏs�`]-����{/U���'�a�q��it�;ڠ+ �i�X˖��Q	:H7SQW�}��X}�њ�'���ϓL�~�Ә�9:-��FkeKs�I�E��R��Գ�y�i��c����{B(ROJa$��<ο�ji�$��0�#��o�����%��"X�8�Hm4�v'�5ch���Jb�D�)S�:�7&�{'YS�hcS��2�*eO_E4ٽ�bY�:{�V���5�V|�c5R�Z�7"es�&� j0kA��2NZ�����)��@�w":�24�zԼ�Z?��!F�"�t�ޓ���F����䂯+�����,�m�|#"�9�v�}��[��Dv"�:��.!��	�O����:h�Jf�y�v�P9nϰE��)��	O<f�	F8}ŁV[Z%�ȳ�4FhTt
�"��~,��x��1�瓦q�u�0��h-��޲M�M�6)!jY5�9%G)�id��[�pguG�r�,i$�����/�:�����o��5���n?g�5\zm�{�L~]�J������q��Ξ���S���Y�~'k^�9p=�,�����,�����w�����}l��Ř���lL��Dƾ����Q	�a�c��DXx����$���V�\���J�`~�;���X׍��T�����	z�R����MlG�l��jQK����@h�<L��	q�JA�G��|w �Z�X��,9��"�aZ�0m�[��ѱ�$|5�Ձr.(Pъ�zb����z
E�ƾ3 �r��F� �/gy������3(+�K��)K�;>�šu�(Vx��ͅ���@Y���T���u�m2ť��n���Ѡޣ��D���I�d�����`�aĠ��W��8Tl���|L
����yV[�;m��~ք̋FPD7�4.���*�A���5Z��5V"'��&��̐�TY�¬�g챴��
��O��r�D���}��	�4�D � _��i�TԆi�t]����g�ޅ�|�3�z����7Cߺ��q}CD�������֟T���~5�c<�G�X��!��U|��H+
tC���? C��8b6ꦄ��S(5��tY�ʆM��b��s��:2'��L:��Ɔq�Z/��h��IY�@H?�fUt{[�:���j�3���~OS����9wE@��~�Ur6�f��*������U7������'̟6&+��=��w��p���SM=P9�1��3�����Z��뫛�{�=�8�X�'
�c�~�ٔo�K��6�Hn�)��B����t���;�z�M,����1C%O����5M�q��Η��<���ή���E53'n#EEf�s�rT�K�Ad <m�S��dN��m�2��Os�$���Hm.�Ul͉̓�/^!T����F�RQڄ�,~�s]��kn];���SHP��Y��/��b�=�e���O�Z"�a���^�7���L��eVC�����!�A�o���]UW,8|�m#W��qĉ��_�vQڮ�M��zg�Lg:;+��;����^�4f0E{+���_m蔖1��툫B��;zZr�S�"��tN3��;�+a!����e��/��uR�2Br�@���E��x�@����c�\NW+��ߛJ n2�L�@
Õ8����ŐS�Mu�������v=@����Xd>�ه{���R��k��8doN$F�/ W����jW�P��:�=T�d�M��?(�[W�)HϢ�����)�!{�� N���X�<j�5�h��{peO��͆E��3Gþ�\�1��-��V�L*�gۂ��>eV`�"�E۲����〨BD��W�H�R�/}q.C����p����X���LK�x2j�B>����Y�DV�dPk�w���k<��C��J���Eu�n=�E��8���(P^��꽈"����I8ݤ[�x背	9��ُ�
�Ԩ/ًT?2� ^_�����1�)�V���ĺJ��E�y#��ΈI��r�$����L�����%��Rw���0G��;|zM�T*���!��M�lc�B��;f������wp�~�׫7�=ݫzr��� KvBY&{�/~���W���<^�T������T��n�2R�J�_�]����5��2�E���[��(��ܷѕ�h"�@�1[�O<�;���h����X=j�hhqNŉ{'Vb� 8-��3{Ũ���];re���Wm��>��x����j+�U��Q�7�J�M�S��ߒ{�y�h�=�{F��ڜ}X��f{�,�����Mh��EfW���:�J���ᐵR�m;(6k3�����4_�]�c�2��x��f3j�1
�-c	�Ƿr�sB�ß6H�ڍH�]b�l��5�����ގ��8|��D�u���!�t�U�|��ﮝrڬ�����)�g��tP�.�ŧ�p���R�g׋x0ץ�ҁ��W^s�\1�V�4�h�B+��E�ߨ{�.�����s�T�s��(���ҜV~�C'��
r�E���l���(�u�`j���&�M7�g[��5�>j"���g`t�~����7)Q�d��8jt�����R����S^@h8D�&�Uu�D'�pQ%6{������4��ۑ����g������ R��&��,&|^+Ob�U�샴�M�����΄3q�A�ykƇ���/G�"4�9�b���4
�J�
�{,܏��N��,Y��%y�f���6X_��"��)�໪��G�ҕ��=���X�wQBX�*��Dh�D�s�J�L��p��c�5�w����W�Q%���H��n f�*o޿(�Z��U��e2��qu��h�7�_��"�|,0���<����E�m�y�'��B-Eϳ�s�R�Iy�(z���)�)�I��/s(���4|�Zz�5��!(��fX�x��V[;f��I=�ԨO�\(>	A��J��2�U������EsV��mbnܕg�Aio�ɺ�w����y�Ƿp �A������QP\�TׯLV*P�\N������ih�1>�A��ܴ�i���G��a���E�n��v�Ka[��>�*�ޏAh�g/C��A��B`N&r\�A���g%���iYi5iŐt4&o�{��ꘔ%��ػ�W�ٽ8�Rz���,���s����*��e��Ȅ��h��c#4?�5���]�*��,�
%A����?����;i=�o8\`���b��
�����Î��{
K)Aw��pLƽ��	[��I��1�vg=��#k\�����ufˢ���>f���ڬx�z�Њ��t[�}���xg�N}o���)0�U��Y)�&��?;�P��5��I�>L�>&\0�����Ҕa��Ͳ�"���K��6~��B���t6�/,8Q�	�����=g;K@I�_n�U��1��25ݍ@+�׎@mT��ʙKW���Gg!'��(ނ5y�[��P:��Y��U�_�l���6�$��lKS(L���lp27⸠�[��MO�`ɧ+\�3�F��`�A��]�b��+y��A:�h���>ff+��ǟ���0,�(��Nfdv�п1Z~������eE���@���λ�Ԣ�}�<���=@e�[���i"���3\Y_ѯs���mp]����N���,��c����o��=��F>poޙI�}s���`.��ы��k%�{��|�P�c�sFI�sz<�ާ��*�Ў�`�[o��>�ۦ����щ�]|$)��T�Pq�G#~�%-����)�X����ٝ�9�����X�+J
ܾ����������qE�"��#˗B#� ��G.3+����X�QJr���h�<y�a��ra�::��Y�K;+R��>Jʻ����S3�Sn,B�"�<un1����`�H$݃jt{��ը�؄���n��i�6�En��Ѻ8w��4kCm8�����=d�K9���M�5UJ�T���}�R�([ER��
vw��S�Z
��M��_(8L�f^hޕŵ��.�P���6�l���_C��b�%�����Ĥ2|EL�o�ӹ3:yV׊P������Ǎߊ��7$d�����h�x[�#@����d�c4�߇�p�̀�h��\���e�(u�d�l��V����2eTQ�Lk���.��aq�Ŭ�a�ǐS�Um���������0�9���Q�>��M#|�+n��Xtf^����UB��"H�@*׮��;��P=��\S����c:����8~�15�1,�?a����k:S�ϗ-5%j6{���e �����o��%%SSRX�.l�ɑ&!x��g��c-����$@g�>����3:B0@@�|>�\��z��P��t����Ǣ] ��m���aM�ب��������N6�;���x�&a�R�ܾfxf��/+'�֘���X��A���	�5wn�%��K螴�ը�*��?�?�H��5�T�>G��b��R�l8��QbN�u���,�"�H�|A}�%���F+P�'nH���~X^������v�� HLy�5��Q�/c�f"^��d�|֦Ɖ�eE�!���6Mw+Yj��W<W��v��?.
0�=Ÿ�}f��6�y4�Lu�Lz���"�e��!�����m�Z��)��$N�=�`���c��Dp�L��1���7P<{��Vl��~S���yŝ�m�i�E�N� ��S[V%mx��/�MUCj��{':՗�& D���&	����ŕ�;_6���<��V5��2	k�nJ7�d�r��V� ���S�)<�����˪�gF�u��u�T����܂mL��dz��N���� ��v�@$�ٷe	ʹ�H��\�g9@T�OA2La�w�Q\�kǨ�Cِ��1G�rԘ
B��ya�4����o�+%WB��p:��C �<�;{�:C���ZeD��{���$F�Şc�%�Z���a*�{i�f��08s�&�,����l�g�}����s_�q���I�o�G���["���J΋>EF�ϋ��;8L��LGI��L�~Ţ-&D{�5�q'D��kr��@�uB�8
Ͷ)�~Z"<Lw6D��[�5{@�R&�� �"��B��9�V蒇���@��4}�(����}��`�#���^��TiE�
��!J� \����ȪbאַT����[I.?I@����c��f�'E'��^��#d1��y�&m��������*��c>#^�3](�ك�A�K�g_�rx�k3�XC��_U�#@�i���k�ƙ���#�$\��C�#܊h�F����%�� 3?�zE���y�G⟆�Z���)�`���~re=���.��e��&��`���2���x��Q��!� �����̠)��i��#T��u�#-	�]��K 
R읺Ui��B�ɐy�2,J���ăOțGF�����XJy<���OS�15�Z	��V�DsB���������V
�-2���M��8i/kJvs"t��!��| ���*�D����}�\� j@�|����d�[���fs�Etъ����@�p����
�qAJ����)i�W��ȿ���o�+�.�Gz�vU8�;��u&�A���gD=)���.7�I	l�cӴ�=S´fO��.6�b�_�P��П����]p�٬�ZL	Lyg
�eѬW�g@�ILs�w$�Px�R���r�a�{�q�xvCLhIw֡����ܘ��-��C	ٗdF�;��wYF�V`�g���I�y�a�w% ��{��
u�l�z+@X�aO��p.f����hFʀ굲"d���E��LW|B���w"~�~c��d����fzy�Tk�4F�y��ݩŚ�"�o FiB�	��e[�c1�D�j%�Ic�k��~f�eY��p_OHjF��&�F�Af�&��5��`���z�M@Z].��Jg�/^<�E�� y��f����c�]r�Ԑ��������4��0�s�'Ҏ���/�}���\�E*� �L�lDna���-���ƃ�'uzzovv�2��к�~O)hr��i�<���a{��<b�3������e������𣁠�Ui�r����I��-��g*���@�ȉ͌rQc�e�cRb��
�����j1��[�4t�S�����`�s�Jea�U��Q}~�g1�a�5�!��a�7��uJo�Y�����+�ƕ��<�DپD~L}�x��ď����	l�!!���ֳ�Q�����[y-�z��͙��՗6�Î�#ˢ�0�RƆJ�;cXB�Z���:���aO%�D���x�� ���W�����������<�m(��u���F.�J<qn�X0�߰.Hkߐ�iO&ApA�C�kNo��/�`��e����O��0�>��L
��׆�#���ѭ�"b=���O���,��Q��F������?�m�#�3�b��@Y$����$��xs�G��n��Y����)\E�Rrr	��@�YJ��?kp���r
�vm�gO�x�祒�J�a���$)ɍX�p������'�I�Z���٠�����v23˅���K���`	��Xm��SF��Wr��ȔSf}Ep��.з)�T˼�P@Q�:J(	m�ս�愎fd-�Cd�O���/P�2����F�<FU�x���T'�@,� e�ySc�j�q�+$��V4'Lm��Tu�y��^�^4��U�}��?Wf�~�j��￷���6I�9)�C'��=�P���g7��wy�������ȵ|�.S([V�lݱ�+��LJ�I����Lbi�=-���P����mM[�čg����VlIOƲz�ߔ��W2' �{.�$��e�I��OP��*�1����"#�� ���k�b]���m\�Ѷ��~Q���&�c�q+����ܮ�=�c G��.Ŀ���4�V�+�X�ΌKĻX��1�y��ur��4��w�j��+��"Lǵ���b�����?P�JeWڣgr�#���{d����W`���,Ղ�\QҘ�ܩ����^ID�n�Ɛ��_�s����$�`����z�6{Rte9H��H2o^hU|&���|$\5����*�V�c�{(�`��f���;r�g9���ɛ�I_���O�P��Ο��g�U��]�W��<NLy�����ݢggo ����~`�َ��
{�[�ʪw���*����D?nz﹝�Bqw
�HZ(r�xhW��y��1�B�#�G{�6�������0�&ݗ�j!�j./���l6;<5;�Y�+w�˝e!�+�p�ܮ#��g�'�t7�L�7�a�x)4B<�7�o��I���ڏ��?)^9�$��<��#bA����[��-�^MVҴ��vM�Xlml�r#�l\[tX��ؒ��\?�����]�mP�o�H��Ä�濸<�����t�~Y�mб/�:������Ė98[����Ж���.��d����z��'7e���"s��n[����1�e%$�#O�H��fI��WQ��8Pѻ������r2�3����S�����N�;  Z�,ʛ�����c��n��!UI�~>�]���[ua(�~�����b�^2��9j�m=�� �?Z@�b���z�%�a�Qt���=��X�6�N�m���G����l]�4�f���f����Lo�����AXESt�Rs �L�J5�U��!���?˛�N�L�V<ͧ�E6���T�T	@E��*���5	%�Na�>GC�z�T�ҶbWqJ��NBq�zs:Lv��%�#��4��
rVy��� ��~w��Ü�(Hڷ��"�x��R}mR&�+�	�s���5��'s;�(�e�J�����#��dM��z��.ɜ���*e���H�D3o�&�yr�,�o�����j�@�N-���I�+�5Hr���J��\�Ly����T~?��&�@:��)��c���.ͥ�1v�)�F�jfl��6Qv��Ꙛk����[�SjY�ω�t��sˈfs�%�lV'�U���W*�Ե/�ZB�No������~\mlr�|�\k���@�4!��5P*��J�M����<�
��[��+����5g�Xg߄������9�x#�;�#��k@�%k4LG��j�����t;�; ͸'�G[���g��R{Lz�
w������ۄ2;;�;������ڥ
7�1up��m��Y�çu�)Ѡ��R��%;��v�y��B!�֕e���E롹F��� (f'k2�l&���	K���h똘�՛�Ke <R<S��ڝ�r;����B�k�jt[�%<7���Q��e�/J��r�"�OH�{iO=���VbL�,��E��#���e{��1(sIa��e�;:�����'�#�dy(�@����a+Y2\防O���p4�p�eB�.#�B�r�f�`$��0�8���Nm"*��&�zͲn�_
_��_{�wo�I=��^�=h����Y�
<��:"�6�/J*�p��<�&�Ș�� �R�x�x}�������9FbS<Y4�|���"=jhT <,"a`�2uT�~��6��Wo�$�
����D8+0~y��Ԗ����Pat���T��+�҃=(?�_±(��y�~�%��� E�$G_��&s�S��Lڡ�R���[%mI�� eKi�>�Y%��
�f�V��RK�c"���
b��A���ϥ)FX.U����Ktx�\�B��Q�x���$QĶ,n��̀�G8�h�I�v=�$
N$�*Y֎E��C�$ �Hg�N�P�6��i�����i1�W����p�P�6���1������8'�}��R�3)�dw��;�V��ql	�5����:")��m�F8U}q�4׷��}|[�n�M	cX�i��fNMț��Ф�.ɡ�p���.s�GC\"Q���P��ci]�]�(��=����L%�t�����rb��Ô���`��� �\(�8�bMƱ�'lno�Ir�
�vF���j�,5�in5Z��{��X����0h�'>;VB=�Y�N�,2e�*I��g��'Ƀ���j.�-�ɑ,A��m�SJ������ ��<�L��|r���d��s|QdO���cH>�q����-� �!;@�7'�׮���GBD$ynR!�� �K��G�@���MèR�I��4?�`����V\�{U����݃�z��/�\tDF��ݜݓ@����@��y�)#�����Y�S��J��o���w�:w�k����fs�}�çM�����A��m/�Z���X9�!�X�$'1b\2�N���.L*Ω��x!�Z`��)�&`4P�wyҺ�u���n������W����⶚ئ2�CuB�|��1M�o� dž� ��ذ6s�"{ٱ<X4�Ӈ%��[��Vg|_A��m�,2_��yhp���iͧ��H�s|���{:s�DGds�߰
��h��W����5��B٭\�q+���8��!��6~�/�Fÿ�R��)��U�KF �:���7��T�DIB$LX����}&��x�����A�ڥ���K�N���ę�&�\��Z���+>�q�f�J��r�i9B��@�����ב \�-�lW����bpq��.�U���~��h��IlSgb�3;��F}`�}:O�8A��Ca������E8'�r�t��,�(89������7AlЖ�*�L$�z5W7)˂,3ke}���vI		̿v݅�ݓB�Y�b����sa�����o�����"o���q�'�
O\lB*Ow�t��ǒm��gq[Է��p�O
�2��ZN+��jOx+���w��+��8����hq��g��w3�{F��0N��}5�B8&�M�g��RXoY*t8�j�
|�)L�����?�����\���ɾ���(Mr!Ǵ�:g�dd�'���t�p}�.�/�2* =S �κ�D��.c�A�B��u��%V*t;a�i������suj����A�'�h�����j��ɚ[�ؿj�~�?��2[�������0y�^�� T�.��쥓"�罱[�� fWKཀྵĨ��;EG!��Z�
��Ŋ�,1�}%2r-r��>W$@X-�^��-�r��dt��hw9�B0����>Qmx>.�Μ-X{�;����#�����oHm �S�A��6d�ӥ|S����д���B�S��bI��r.�=�,Z�v�(`�~�������`�~��(���[*/x��=��'��6�(��땠Eh�x�'�=�Wj�L"L���*;q#��b���fk�aw�m��
�ତ�ç�Q��0��1I�+ �}�� �����旅)�6�^7U���wh5X\iAe��"�[d?A��?n�S���(^)�Pk�)������P���_E3m�e�*6�4����$�����R.+t�\�I���[J�>H�m�'q�OvZ� �um��2��f�\G���!^@���W�����F��Qt���Np`zr�c�l��n��Aj(��]+H�S�q�j�Mã��Y�x�Rܣg�mz�� ���b��nQ�����Dpb�
"��v�V2�-���>�����E�����WQHwH���{��Ꟈ���X��k#�����<'����nS>���G�! SNdl{p(����U~+�_t����
�VVR�~� ET�5�!h���$!��fO����'/`��^Ƴ�������@��s�F"4���蠫)�J�a�����Qǈ>���r��<��,0�Cco�@��֝)U��������7ɛ[�QoćVb|�*���D�\d����v~��+�pI�/9������n�����$�'7u���S�ih,�x���1�Mݍ���n�ح�hT�3�=+�"\����\d�E�;�	�]LX���[.5b7�=+lN�?d1�ˏբ�N������'i��1���=�C��0*u��7#|���tǌ�>ꇂ��V����w���n��/md�?���j>�!48ѵ��]�pf��aQ����!�S�ڭn�m?0�6wM#}|�0�/hXkaQr�����.�q����'��F��W�c�4�Fi�ĞJd4�m�42�H�zڧ�м�_��&�P/1�����O?��ik5jf�[?�spҨ��w-1����{C 
��6�#׆�#���/�gryx|�c�e6��Ӹ�ҏ�{���Q��n�%4�S_;��X��w��Xur��	=d|�� �,�:c=��$��i��Nm��9ӝ)��8�-�ƟDA�~ ��rݍ�-��y��3w��v�}�D��W���� �
�t1T���rڇeS�ߦ�GJ�%��,B��!�8O�Ww/�X�����Z���R�Mwum< ���֙�-�rL���<A|ʹ���~�-�A���"�n�!�Tm�!�����&��Y?��P2Zhdܲ��[CɓS��eMm�%��}Mٮ�zsYGL�w}�=(�0��|tu	����r��Ωߟ�F�ѡ�T�
�)��?����_'<�kDd����8�O�Z��w&�^Q���\�z�.�m�JA�[X��V"\neغr����;Ѱt��փI]��ɻ���ר;;�o������`��u!m\�9��6;{&��h�Sq��u�cT���4�Ig2��x�b+�l��R��ͣu��[��e�����	�w8|�5%��G�!
�JSNːQ1��9�夻Y�
+��2����'vo��u�����
�GaX���<UP�QW� g�`o2��QYG9uE�/�I�z9��u��p��>�X�����ǿ$�GBW���(Co�?��4<���:�6|x���� ���	I;�T����E�C]ae�	q��2� �:M��	b��c�ȟ���@�8�'w��q����{PFT����`���1���Z��9ϗ�; $3ir�!�M�4�92�wƊX-�]���k��u��a���-l-�����}qx)~�W�0�v�x�k2�0(��Rr��q�m�C�8Q�~;?g���,��LH�p�-�G�H#܌M���I;{����~|�Ro��b��QW�g��x��f��Vt�3�n���Ө��:\��*(=*�0��hc��F�Q��JN�|��?��ȉ{�8k]@sL�9��H.�E�#" �T�l2��e�[�	��<��	���¸������U��g�>���8*��\�J�<����eb�ûĪ�(�L�-�,�x8�I��-ߗ���!3��|�f�r��� �n��-����tS
 '�*؃�;|��}�i��8!BcjxO��RKv�a	lǺ�ʪZ��l��'�}���3{Ca���CW�<�D��Gc�@�vW0������=tJ
^d`��h����d�Rܽ��X�W���c�FId,��+d[@H�,���h�6)����T��ڴ�,�$�m�諆:��4���R�m�
��l���q�*t�&��-�kf��G�3���\����!Z�ͱ�����^Mr�����N��5�� WTr)��^V@CZk�0�Ѯ��ѻ	t�综�����=-8�{Ho���O���ъ����m�V�Or��
*�YxL� '��.�.-� �Y��յ�,�2i��1�!���WF���F�;����6�dxkm�x.�m�;��c�WT�$F�y�Ao8Д���07T�;�{R��J6㤳	vQ#�:�by��q	|�(鈒,����u��&ܠ�b��[���Jnz�1k��R�y���շ����z�f��!�IQ/T��w��`��Ӏ]�i8[�-w��FVF��H�Y�#�	�a_^��� ��Fҗ ��esvƽ��ͪ8�S��<�Be���z �0�����&�#�TBU�h�m\���3�$�9�O���y���d�R�<"�F�:���$)�I���30����Ru]�U��[��X�`ݩE�����S-�5��$m�4���M-�>ѷ��Kf��Y�Je&�z.�\M�����v�I �YЛ��=N���Ŷ���\�$О��_�_�H�Xv��C����ɰ]�r���J0zp-.��M��v��
>�� �o4fٶc�G`��h�v&�$u���)h�����r�R����D徹���X�:e���,��m@p�i߳���g*\Q'�6�Y�<���=����WR�ꥷ �],�u<	�(��BxB~�L�&��՗u�ޏ���w�ָʪ�
�	�)��Va5������ݧQ��* ���xԢu>���$�uZ"[h��J��w`�£����y8��=q�V��#玾!�qs����dO�<�"$�4t�s5c�]·�������jh�p�),mЮVL�z!�Vf�5�6�Q�=����z����B���Sv�9K�V
5:���"�\�5��2u��j}d�Ԭ��q�C�zYT<�W�U����M�*����f���C����l���KB�h�	q���>�'f�ã��G|��������K���%s��2���2�6dG�M���t�aC���&��z����q]�ܜ�x �����.�h@mK��4�:n ��zYj����nB���?+b�Fp}6�3�^��~���5��:6�N����6����)�h��YZ�����,�*�$���0��&LRo�2c�uD�Nu���F�Q]�౽=�d�_du��I�?iXć����6�g��u*<ld�Y�/��XB����@ҍ��,Y_�lA���	D�&���-N�x�M�'�$�Z�ȍ��j�Ӻw:��,s5`��R��t��)�n|�_���%��8^G�v����ɋ���ɬ"s��2�5W�.�{^+I�k�i�����}��{8�U����?�,YD.��b����9K�[b'U��A�Q��&P��4�DCܵͲ�֝�L�";�� k¾˟��X���Eö�`�#��^��_t�~��m7L�>�'Ɍ��,2��;�K�o<q�(�����=���wĪӂ�,ھ=s�ȓ��av-c�y�Y�9'��2:4���4�J���'_]͸>p�̖�����DR���Y��S{܄q�Edhe��*gC�z��7�`�<�K�`.v0n팟�tg�Q����>_9Z�C�;�>E�R��{RiE��m@�4>�B�f��ᝨH��m	i�av��R�Hˢ�j��*b
��yH�6Y����014��<C�t�TJM|W		�������ܺ�p�
1�Bq��	Tu������8�DN������qB��_�.���G��iNimS��fT��wLݝ�����DԮ�����}�Lzj��0�Y����\H���3��6�z��)��i�����P�E��I�`�D���H�6�H�'c}�_E�D�AܴӘ�ɏ�!�wi�.��t �W�F�v��"�� ���w��W|�]~�]=�>�zmV���o��j�4��\���O2�d&�8-Rڨd�� wty��WJD�2phO��4��UpY?'ׇ�y'%O�P�Q�S��	�E��՜������,�c�:,�Dd��\�F�Nl'o���F��W�q�{�7je!���5V�	٪s\�ch��d ���(�vqA]l��E�s{AVo� �� �j)S��̐&�-�������C�޴TS��t�^��D����G��qZsy$�N��g��`��f�wu�䗾���N���Gubf���7�OȐ�?p
��e��ȨR�FOu����Y~5���3��.
����j�����Bl�j�< ��P��(��\HM�];l Ӧ{�*g]��^Q$^3�OS�����fD�0��w�R��3Kx�N��Kڅ��6��U���/��l��)����$(wY�Y���3�>ݏ�I�s��s���x�
�l3��2�ؘ�+�;�6¼�������_�[}��ӏ���r�j���Q��r |�W;A�k2e�Qj�j�ŝ�-���D�B��7P��[�v7Pli��x�6�5�^��R��:�<p�&{�0�?Bk��s�$@7n��"� ��3�����h�f����\��&��4��W�Q���� �[;�aqD#c���nkW4췭%��!J5�v�Af�b/,��b�9!���8�s��š���v"�����P�Z0�����ɊE%T}{�J�ۊEؖ��&"8�O)u0��������A0k����Q~ZHpn1��?t����q|��g���'�o��x
o������x�:�%�Fa�8O axwpN�<%�6�n�ԡH�*M��W� }i��ѱ2�g�f^9�}+��cL1�sw��ý˒�FrD�Kv�B�.l �_�.�P�&,�YUq��=z7�A!'�8x���^�s�$i�2/��R+뗫M��l3`�;O��D\A��� Z�C��3Di��U��0ep�����z��*�~l�-,u�)s:��F��@�s�_�A�3x�>#'�`sb/�a�[̢Q����ِ���5A����0s�E{�1�Յ����-�\İM�YJ�|��`�pE�ޛlk����HU���I�F��2�ϜJ�\g-��5�)�Cb�L�|�)3N�,���}�������MEEOOQq�XʚZg��q�W���ڮ�~j��AG��Y�!��;0w�t���H~� ��� �'=��	�@�)3�x|q����?�<R��*Y�NY�q�՗�1N��n�ɝ�N<]p��9�trܚ,�����#�����ll1`_,OA�	�+���ק:Bh����E|� �1h��(o��?���ی$�Шx���.�T�u=�����&�~Y�|��=��K�K�E�����M	%gZ�a���R��p?��U����-kE֊�]����ίf� ��}�%��yޤ6����ja�j�>6�.i�!��:`�1��l�l��Pu#A]��/'Yj��SV�~iW��"u(�4��w�;�K��|9�^˦Cm� |P����ךNn
R��l֊8Fl\�,�W@�G ����/�R��T� �<��τ�[G��na�S(Y�׮2���~,?+_�2)W�U�� ՟0q]/>�:M�{[d��0g.{Uy�x��T��%;��iH�%(`L"���,�W߽���B|o���Kv����.��r�!~`�A<�]$��Z���z�r�H�����Aјg���<���0��6���[6AI�
�Q��F	;���	��4�ں�ñ_�u�C�?A��C/'Lf	H�x��B�eTG���i��H���ﴁ`/���������E��?<6�  �,]|;.$��W�L��S���Ј�t�>��&���p�j��.Y�A
-�	����?�C��ı�/�@�=S�B���lC���q�1�����1M(N��ke�Ю*�@Td��s���d=�%�#Z����4��ꉷ��)�*��rƚ��[�}Cg����yߦ������O�R:	BO6�򠨪����u�!v�I�\P���S����<���e{� ��\�q�1}�žC�5�y���Orw&�X�����b�;p��V�(.r�����/;ҿo�����P ��y�jLeLA� g/s�d��+���S�R���K��J�^f�M&�(���6��'VK>��N��������q��X̙�`�)�шwxZp{DB�)�$6���n�F?��s�	?q<FJ��a���u���'�f�%щV*��Y�e f�h���`@4�)��/��\��
S�ȝ ��EB�#)QG���
ˡt�%����Ww�(OX���a�e�l�7���I`��SL���:"�H�K1y�)���\�
�q�Bw9�p~�:��
�NA�jv���2}��'�T��vn�0�J�U��%H�������,�E�m���ׯ8��`��e,m#}���6ܒ����W��m'K����R)g�E��~����
n��ٜk}	$�b2�j�4��;�\5������$��b^�[IfʽӚ�P��)���	�ȶ#I��]�iS���=�V��=$j���z>N�޵�^;k������TZ���9Ն��V�׀��}�D���&��wu���}�Y��uۆ�8)i�"�Kڍ�'_����3�0�&W���c8�~��љ� ~�j�MEs�C"���vi'*�q4oP�r�a�!���&�z���M�:g�R:~�T��0eT3?�G��NI�	�ߪo�ţ�ycZ���ۿ��5�m;���9<&�jɦU5�����2j/~; �$�Qΐ5\¨�L��פn+��CVm�Bں��ԝt�T��d��z�W�;3��{�tD�� 1M囑�\�)鍊�e;��Ň�lހ5�鰵�x�d
�����S��e[�G��oT:�Rv��]!��!9��s�
M
��Ct�j�#���4k/�*hrdn��1�	{ZƊC�j�hcMl,T5��-imf���g�C�u�\f����Q�
e���t�X~����휰�O\7<�֠����]v7)[:��q�+�g����7q���ʛlm�����@Q!�X��[����J�!��0OuaϹYأ1�C����Ƽ��,��	Y
��y�Lt*���h���`�pQ�7�¢K'���E����,��=����g�B�s�ؘ����$������h�)�3K~+�٩$�gs�5�$;M9��h����!V�V[�Y�&5�c���uݜ���!�_X��M�Z�v�|�RE{ ��6��~��h^�يe�6iHp�4B��V���7�`���=G���i7����%z��v���~����YW��fH�	fݭ2O{	#n�1���=e���bT�#"��'���b#�ڡw���Q���v���qX�u�����o®��̩�#M���Th2��K�j���H�:D���C�����5��f|��5�b��N�\\'I\���;�?�Fo�Q��.�6�YS�,����ه��8s~V/5c1�FN!�]�,~|Rh����$�lv��8�E����-�����D�s�ǔg�������X��J�����S_Yՠ�zP]a!�rů2�y����x^��9�����*`e�"�p9E��%�&�Fhc�q�]�nN<��,����pjz|2�D_�h��v��n3Ʀ�=1���)�$����'�H�2�g�CʦX�M-�YaA��	�N����>��$�th�M��jbi�������u���Լ�m4�D.Y}®<8��1'������[�9(��ŭ�2*�]�'e1�$�2��m/����qO�&��0|D�����FP�����/����&�.�ʤ��26H��+�v��1/��)0��%�v�/,�Mhsһ�񶤽"&�&G�Q
F28�9��O����pq����F�AJ��r�y��6����.����UW.d�9ˁ����������_D(W�F��RN�B�}��蠿���+�ɎF��0j��8��<M���H���k��6���X����
ԡ��n�r�QL�_��,3�~��ӿv�Y9�3�ܦkp�򘣖��	r��0kFbƀ���	�>��7�6�1�N�&~�Dv���c�<o�����F��
l�!$��+��$�	��#�f��A_,��q�t40�q�^��; ����S�����?���K�:�%�
�e���ذ��c���(�a0�x�k^�1�j}�]���r������v�&f\ �M����d�͵a��pA���W�瓧���]`��+?c��[���i�
�����6It�	�����uҀ��Qo'ĩ3MAOC7��C�ы�U�k��G:Yw%3�Ub���	�)ؕ��"���ۺɩ�6l�p��1T&ŀ=|�t���g�t�^EюG^�j�Oz��0�^
H�K���%Ҋ=*��E:&n
cї����<��1:�Q>|FP�NZ�"V���}{�p����IV�z�򀮜h��z�݈Vݡ���P̓FOb���q��)��Z��E8�L����.*_��S���qs�C��
6!|�M��OGG��/��L��V_�\�G�W>���#�",���_v�D�B<Չ��ī�.�Z��K/K�s�r4�*?^+�}C;H3Ik����6�9�,�4i���e�6|,�	��1��� Q�۳V�AM6^�[�������F oqE̦u�$�����"5��x���C�܌gf���t8�rC�r��o5Ǭ=��n-?t�O'����:��^Y�\0g����j�u|��P�ra�����"d5-��7��� ��.w[y�
)|_��̌|֖;��A�~@���ix ��0��Uj��H��5 ����Q�W��;�=	S_�I��sg�&�"�1t6��K���5s&ܡ���sC��������'��"�@�����} ����7@A��4�M$�ǥ��]~�-̫�	�7����A�e���?���]�a��N� ����p��W�c�Wюv�-�#��Q�%����W$��uo�o^�M�5��̕�����{HҤ_'�T�(Ҕ�q���S�ҨQK?I*y"NzS"��=z��{�bDS'�$�Sy���$$�%)�P�N]�'Hd�^	G�5��� s��ހ�c������PO����=�F�ܣ�&��-��}6�5z��U{[�ԍ �r����s�Lo}�+��U�' �T.Bc;i�*J���?��hW�G�jG^^�-��I��Zد�+��bӁŮ��O����%7�b(��(V�Ąh��	��a�?� O��1	�Y;��=�!1Dż�C���,ջ!1��h�[���k���&%��޷݉M�C-81*��k	"��p��j�qw<Jxw`_
#ui�I�QȮl�d�c�2F�W����"�s^��9��ӛi��T� �r�ĶV�ַr�l��+�5��Մ��l��r<TPI}wכ�C/)}�y����օ���Ck����"#���*�B.�C�{`HЏl@��,��D%(���c���2ZIU<��O �U�B�#�����\�.:}���V���)���3��Bv�	���%H��<�h�-���!���x�tdFIa��ʣ�B$��;�A?p�BX�ƾ	i򾆠U�Pr��4Yoi1;��ሜ�ºW��>�'�[�=ԃ��Њ"v�� 5S@#D�n@��٘���M�:)/����̚�C��:'��X{|{���Wt,+��%$���Q��|b�ϧ�k;�F<�B�g����B�av\̙��9�����7����M9��-	�[*���@�t
�I��;����V ���)��C���Dg�,<��+P�q�#f�޺\��>	ۉ���bHe�i�$�Jh�&��v�EO�U��p3���7�A��3K���q:������l^��ͺ��xm�ݯ������E��)�#d9���]�y�u/q�B�HS`���Nh�0��L�c�1x&��A��V��R���ف(J'�>q�n$s�)J�EA��)���h^B����y������$��z�JHR�+Zݓ/�Gе~�ca�W4��t-I�����v�K���:�|EJ +�r{�¿���9ư��x�TQ�8�ܿVO��N(�Nc:7��0����F<KM�Տ��x�Z�NU�)z�]}e��!$M|U-�la�5����� F�Sb��n����|���{[a��V��&i�	��������9^�I��.];���Τ�dR�`~�bA���9��_� ���Uk/~Y����8�@�LW(%6]��ǭ�A��3��i�������v-�Kދ��kٯ�S�Ӛ'�|H%�#�����)�p
W"{�B��D�[K��/P�F�_�p�XXZk���X�s5k��ֈ�G���
�_��p-A�I���$t�hZw4t�c�=�u�1��DU�^Ml�O	C��i�7q�߇���*9�j��7��[��>^�DE�ón<��*�(� {�*=������TUޖ��`�3t�,�*a �;���Q<oY/Q�;w0�1�*� ��-z�а0\�iP�2��p(�Ģ�pAR@�T��a/l�z̟�h�u�b�L"-]?����X�`��_����jZ�1�� �����VV��/u/�������-6 �j����E��Lօ��U���7"m�p�3\4��N3�q���EM��>!ݽ���\�P
_1ؔ�5<�����ڈ]��~�w����$a.X�J�^����%�UL�.���K�l�S�L�͊H<�D��x�|UDt�̇�1�����*gj�Ň{����W��RP�d��>a�'�'��Cԉ��@+��jC����R�M@b��w���g`�� �ȗ�|��Xp���lt}���z���Te������<�o�����>���'�L�RF�ҥ�X��6�<l6��W�t>��!�bކ��,����J'&��up���K�`ÿ�	e�8�����{O��r�aB�I��zS�r0@p��ؓ�_����9ƥi>@��iζy��+G��;߼��]OA2�?Y�/u��ӛ`·�1p�i� E�w����%�kaxF�RW!�k���}d�O�gIh�{�9ωw��أOڔ�U��P��S�q�W�-VN�@�������/E�q���XV�5<b�;n�e��Y�Ӥ
��<�]�@�R,�oϥ����	~��5�m=7��އ��ٺ[�m����F=´��L�+�#7�`�{�p�n�1������}�$Te��d��l�	����l����8=8~t B��䙒���y4��vv�5qQ�p��O?C�\��V�$	���5�,r���T_ 09B'�-�Ƕ,���D�)7��'�L��1��@������eT�;���Qei��*ᦝ� yR���,𻴪�F�%��-�A��kz�UXq�
ey@=�(�"M#Ix��h]Sq���_H����=�Q(gE4 ���Iqdc� ئ�/���i��YZ����U�U}BXv���x��5G]kO�h]:��c���SQ1*fN����Z�����ɇ��*��	a�^��r���ъ�o�� �6��NФ�飍y����1s��>X�Y�2#�@Շ1x|�A1�-M�_%�)qQ�8�fu�ي�;�G��yO�.Sis
���y_LWn��7�!f��ͣ�?���XV�$R��(Zn�s_�a=�e�����RG�������5��_�����Qy�-F�5v_��x w�q�}�<-j�<�����JL���I��w��XN�n���a�_�d���̬��q��Xo����f���/���r,���y��&6UGE��.���	�yM�(��li�ܑa�Lʏ뗛���Cl6 �/�~ڶR�]��;�;��-�p�n󔸐vn.��Kǎ��;�ʸ5Y��rH��q������6��Oڂ�4�iy�D?GӪ���ݵ�H�CFgDs���u��k ���/����4���7��W��&}I�\����
:z��t��@�(J����2������/7r�)��(Y��`����D��f����5tM�-.6��"��m���]�,�W��~�M	���n�4"�]���U[�Ȯ�_�iX�TҜ�͹9Đ���R.�Ԗ��1����7N�hbg����1����Iכ|TT�&|T����F@%�Y�o�T��.�9�� �9.��,.��Lp4ykQ�HTL�U�"��5aT3B�(�_�ؓ�x~�x-����+��ݠF�7�h�'�2�U������,�L?�
TM�/w���0��G�Q�R(/ա��F�����N�,�Pu�<�Q���Z��<��+wK(��^w0��9B�Wi���<�A9���|��f��5H�F�/�M���;U��k2�q�9���h0JTq��a�]�$�"���i�՝��Y�zc	��U�3�-~��U)갥w�rg��9�K�o��z����
KbV��a���?梏/�zn�oX��i4_�FLv�R�aPʤ���pN�l�"(�cv�UMbP�Qm��X�s��:r!)����͘��7kK���_-)�I�e��W;�%�!Z+���1k8!8P>�W�h�w�{>�̶:��p�zk�A����wZe�0R+��h��Dp����B?{��x�9B��[�dB|]��ɬ!��\�#*n�X�̻:ޞ� s`�?a�3�ڄ�؊6�FT,���g>Ye�hk�[8�;͑�n� ��9*�ڨ�zv��N�,R�q�9(�
Ӽ^243�*tRR��4 �%t gbM)���fu��&��ݜ��9�7
��m��Y�ktp����OO(��3��=L7m��dg�����ݵEu4%a}��7�J|��o_L����55M�C�j(	3�s��6�%z��c�6. HQ_s��ƏM$�wY��>�>Q�p%	���@�� /Ѭ�N?ݮ�G���A�禘�9��ۯ�����ǖ��ðbC,9��{\gW�diʇ��cQp�F��e���:��>�#�.�R)<�d.�3�	��g�������s���Zַm��Q��vsF% #�<Cg|�p����:�Uج��(~����U��D=ܠ��< G���5�_�����
��5�|26�ҹ֗��]Y+����"Hv#����N��a0�����^69�{����ݬ������μ���L��b�^��i�f��B�;w+w���	�S��ƻ�ߌ�q��dG�T�G� �����L�r��uH��%#������ac�Ø?�6���[��/q\�"v�C�`	�S�H���%g5� _hї��L0+W& ޕθ�e�x�j�Kx �u��r4�o%<#�'�R���F(�����7鎿�\�~s�ְ/}� QO�����hU�����h�HF3�&q �@6��K��P9A���L����T=��ٲ��)�N"�`��x�0X?�W�����!�;s߳2��㳾� >�g��O�Ţi�q�6� �hx�﨧\�as��z���_>�����HS+�,'<���hI��3>m�b#Ъ$aOX��������G�:�Y�)R�^x�1vT9�/��UJ�Lgh� �����c&k��9�ai?�F��1��"��u���WΝt��v���D�̹��{x$awP��%�H6��jZ��ކٽB1�����x�:�u3�^�|_*�HE����}נb���ی�n�7�_�[��D^���� Q�@�//G�R����@x���0^g���l��ߏ1=�kz1��*�4�6M�R��T/��h�U'lx���A>�����<Vw>'aP�d�8�/�0Q/�����/���3���;*�8y&5�6��E}'�΢��:B�R�`��cݰ'2����q14�w1G�W��W�X��G�}��Z�u��k i���6��Ŵ(\���}�z�TPR����G;�<
���Sޜpr�ȯ����;�k,�	8�3d�g�y����>y5�9ە�����_�d�Q��R�<���Ր8�Yt��8G=US�	e�I�#�0W\�-'�\���+��t���?x�G��6��OC!��g���ͨ�4��-��Ǔ��6?������+i��5��"ZӪ��7�y��j���:��O��_I�*W���ysK\�S�M�_������m�b�:k������l_���nN�w��.[�Mx|��Ab�)�2�@S�E	$j�~�|�l���I�Z�ۢ�<)bD���+u���n��F�	V�T�"bդ��7O,8�cdueX�PD),�:��k�YW����\�ܒ��'3Q$B%v(�w&�Q%�()P5��16h �%8m17�}�OCB�Ƥ�7
{�FM"?���N������7FpS��G�Ռ?��5��x|#NS=X8��褦W������~_j����4Ǆ5/�3�3yQ��Ԙ$vk�<�l4E~)ڳ�SZ��k����H���-�Y��k�y�X6�J^,1���U��P�!?�N�R�QY���!��B,O�v��%����>�}�W;��&�鯒+ڜ}L����	�D��Ȓ%ڇ���4��*p�6b4����i�&�)D������ٷZ^� �� VF2�M<�JB�'�k�̌�����a_�h͜#��yGҤB�L_A��ļ&Tq\�q���`J�
?���I����"a�Կ/�Sh�;�*�\&�+~�,ls޴z�u2z��d�G�̼���*�{��1�ܝ�BGbb��:V?��L"��'�i���?�$��0��((8��i�p���@����N;�Ϲrn�6\�CQa��l��&�}�+k�������./��>���'�P�����q�RbL�1��t�\��]�j:�M���?��a3o�t)��F�-�����mT%wE`%�jI.�����f�'N9v��<Tۓ���cD*���f���I�0mU���2ٴ��ׁ�\�ӗpI��}�Z��>/�I;���������v_�^�-&��ෙ��
�ف! M�,-���3!
Aτlu/B48�zW�֊��J�C�i�Q��2s]�LQ�'�f^�P�V@�u�H/n�FZ�긒���s*'���s��
!�}���r�Pp��n��4�Ғ�8�A�21�^f&��ʜ�,N���c���H�}��wl�.����LJ��
���=٩6zB�h�͏x@�{B�ǾA�,�����Y�lL:I��$	���X��.9Oڷr�6-��7b O����sf�^��{T䖻Db�j*�r�Bp���VW!bl1k������͇�G��F�ܺ'֫�r���;Sp��.�H��&QĢg�H#��R��Z
�.��
!e7�hCч�4�`���0;�Y}��J�s�a�׷|u�-E.Hb���}�9�)���m���{+��0$������Vb;�Lm��b�0�r}Q��.2��{TB�II~�&V~윁���J��vAB�>q�OM�}lc�{]��hrA�8B�8?V���S�c~�p�q��J�xB6(��Z]/ADړ���a^;�ލ����[j/��C���D�G�]?�g�P����>XXP�F���(%>��el��$��V��k��N�g�Z��lp�N����뜼��Kr��E���ޯkb0��gApÚ.����PR`k�VC&�m�V�~����y6�����ɍ�70$�S�O�U�Uv$t��A|��\j����8�A|.|�����dtʊ
�T�h����d#�d��I��G��/Y;�k�}�B�U���a���0�O�����sQ�Semz-��=��o��k.?�����'�|�����,|���L�O���8�+�[�n���5�b�-���
Ý_��Wf��}gU"����&n͟�ڏ	��\l�C�]߈����΁^NT��{3�݆��bq�����w�Ϛ�����o/�L�ʊ\oA��%��C�$���/�o�@���l0�AeQ��K-�SJ�گ]�#�l�h��=��jyi�E����pj3�Ca����Hq�t[}��7�G��s�m(�o�߻x  �\�<���H:h︡ߪG�W��d�&.M�h�n\a�;t�E!����7 �ڃ"蟖���<R��h��v��b�'()��'�� l�j���M1�!�DxŴ\��P��nP���tm�!�C���NR��"A�F�W֏_6�"JǱ��M��%Ë|��C�l�#�Wh��o��jޖU�&��S�.-��� Z�� �R:��%J�Tgx1ޣ���m�Һ��p�(U�!�-2�S�Aet��4Fjyb:H��Ϡ/�e����
1�i�?����� ��o�*Ξ>�*+oA/��[��``�ٓ�%�3�o�wf��&�0v� y�|�Ӡ��,	��-�R�˩��w�(�K]y�/��T�,��~HSi*!�T�X�2i�&��I����?J ��F�<����:KJ���$%zl��o��vZ\i��^<[��#&1!�]퍤��C���!/k�([�3y~�W������t�&N]�M�$+gƎ��0Po՛��x��I(�n�b��g~�^�u�?� �5H�{w΃@8�m4a?�I��"��%f�����)ކH�������P���t� �����n�S.�V��x��3����'���������:fw=Y�f�&*ԑ����7��ݞj�d2�m�'G���a�@�W�,�^J}��]��tO��5Ʊ��V�E���#��@T�f�|c+5�?p=3��[=P ���t�����]�Y{�ɜ�X����)m��Ϗq/A[S�I��`�,�g�yj���@47HZ]�'�=-�
�d���u��8`���w�z��:}O9N���m9kh�o����.f��C��J$?`�4�I�_��LSx
�R0ly�|�#��k`n�dn'�O�J�8�a;��ԭ߿���4PAB_�!<;��M�sz�6�u�������&�Ư���6�#o0��uR��Rȷ�&�m7A�M��VW�ƣh���\�H�1GWr��i�z�� �ЭB���ۘ�{�XHтʍ�S� ��xP��p��	��h�Osx�6�ţ1�3����=�[��
ƽ���"��;�
ePYI��s  ���6.����3&��fq�i����L�߂����,���7�Go\U��O����bz3�9觰�`*������Hȓ��h����?^�;ixB�%wo�o;^u����L��0�0�P�p$�N�n�K`T;]}@�+�]�C�.�;��2�A���]��TL����N��ͷ.H�=�r�g����7+
��i�\��;{-�X�.Q������o#�=����3��W������2Q���`���iaIb����z���ϟ���9�^D���Y���25���FZD����`���VP*~��z�Ө~B��sJS����ůǣz�Sk'_�"I�C!�J��|�pR��[���xv-g�J����o�
8�'N�b�ڵX�J�-?f��%&^�����*x?��N��z��c������"���(Q������M�3��h���F��o�S�~��wt=�N��O���?�=]ϩ�����;���` �V�(R�!��`H�Vq�bA�N�&L�PV�G���ٳ*��*�L�à�B�X1�.@{3����P
�*+X�5��6*x�{U�yd��{�����~]��Y��h>;����I�7�Ӷt�s�'m���0�G"涉%���|�ܩG�|0K,l�4�žL|w���|1��iD���;%\�L�ʅON����Q���z�J@��ie6 ׍�Ŭ �������׺�c�Zf����h���s���B��	���)��v[�,�@$����[ǈAa�A��Ca��:���祙jz_����k�sA�ߍk�M�<y�0��Ͼ�^ҟp�B��0��a�ݰ�FKJ��@��T�W8�`j��N_d���κ���t��p:wD�oޞ�U�A?n�j~���� ?��R����;|~���� �r2���`L���/Ou����h�d�K�Sr�Wᖽ�|9=+$F��Ć7]K����mb׽�+~o<��_C*38l�lm?eΝ㠾t"�^O�Ѧ�����wΠ�L)I9ݜ)�%	N362�]`�W�������0����}w�խv�!��;�M��hV�C�����wH&�EX��Yƒq���|�a����GmMyUY��$�!Z�����}���9�Țz���ÞJO����{������P�^s	�+���g��ո)>!�׃�g+�4���)f?��b#9�;���Y!pM^4���� �3
q�v�YQ�19���$����\��ZG��<}ƞ���}��I(�*�����<���u�$�	���|� R-����%`��xۛ�C��+���ǟ���m��h�|"�.w5��^lFAY�@�_�Xm�jѿ���\�"��Go��/��ĥenc	��U7�ס�a��x��+���F�J9����n��v�"8����+���𯝇c��(pͰ^�&�-�㌣ �p3Xc�U� P�ͫ�z�a��1�{%',��}�_U���zd���c|.B���� OTU���;��|X�A���F��E+�%�ԡ!Z6����qwo�?���ͼ� �>|Sb8^*8	�(8��'!�
3o6V�
w-�!��+"?�(�`�dg�h��6�&sb�uw�D��D4��S"��8�϶ȻN��]8C��7O�w4#g!7j^��\��dz�)����n�0D���+�eb;{Y��8����\������$p��x�k�ǡu�/� q��w�����-!��$��J��a��!�����Z�/���I��n�;���:����)�s�r��*���^�,�Hg�+��D}���*ե�:��/������h���b�4���ι<�T[
[��������P�>�d��=��xoBƇ�
a��<����\`��\�Ժ���ı$���d3�4ѓU�x<�:����SѢ�G�[m�~W�c�EST����N�&�y�<8�ӫ٭�[�m�e�%n����#�&��@L�����A�l��ҙ�-���_{v�%��E�e�=E#�����&��Q��Qd�ԛ9�Q�����~��$���f��?�y#p��ͫ�<�w����o�� ߕ�B�fW��tOz���C��*��or~�w�u�{W���(�Q��x���G~� «�s�>��7g�ވ��^�j�I�����1*ʖ8���Fp�\����b7�c8���]
����M���������W@�"�i�Yݍ�_"� >�����^�V
U��[A46)Ɍ'd���5��J��e�»P*&)���Zy�9}������"�r�q�s㊌����@#h`��[�3��7,@�'M���D�,Vۘ�,#3Y�	���V2N��c:�ѧ4�"AN"m&�!]��I���z��gPc�P�&!�^�7�bN���5�z������ą3�Í�	�Rm�:�F�[��XmVƩ��'�B�����'_zz؞k���.�3Y��$�l-p��"K��	�*�5oD2�<۷�&W%x�����3��M�U��H�\�ۏN]ܛw��� �@�ͼ����
�vv�s��U���f>6w��ԫU�	N�K��)�M���զ%��[U�*�s���wG���\�ه��P���L��Ab�Z0x7H��h��5;�l����[8�1>�	��m���R`��W:�#�Ѡ��B��h9���lお��N�Mb:^/Q'=~+�iv�k�_��ج��lD������-D�p;q�d�qF��1���;n�~b�>\xY��ZD���Za��}/@|�?UYG�+����z����@b3 ���4��
��(]`ds5"�Ё�ל.k�Զ���1�H�ON�E�tT��ry��C��쉴���w��Y7�do�y�q>M���_�q�M��n1sI�:(;*!�b9�hgL��!^����t�]���x��~/@m�(��q?��HY�n`T󨕕��R|��n���ǥ������Q��K��ȁ�c��O� �_���˗?�t�X)5��i<���u�?Qz��������\�4�t�=�@�Hu��v�=r�3�~Ǳf�{#'�K�C6�G�>�=F;l��6�?'/�E�q|LrS\�i���&��z���X᱂	po�o� �X�2��T2}���P�B as0 6T�%nǱ]� :��/0�*y8��5-�ˈ�<u�ٿgҴ;��je�v8�n�!�m��ٱ�,ݽ���d�ށ��r�T�Cf�Nj��$���%�ַ�_��:�ӗ/\�&Xւ��5;iZ�<�!����Kp4�x[6S�S=R@W�b��(v�@��Ȳm�[��H�Rj��%Ay,qO�!�L�ђ���3��(JTpD.��� �(����ZӜc;6|0V�9Aգ�5x.z�9�0F�pZ&����W�`9��!@�F�z�?v����X���jQu�yc\C�9N�*	��8�yF I���m�:�1BNe�ߑ�t�D�	_��h43�^J���.GM�3O	)6�`C�a�g2�L��������X��j�^vs�Ŝ,�ȗ6W�;:M�+=n�!\���s]����o9}��`�XYr҅L��&���*�hV �2^����L���B.㾶��jD5�K^O:]��#��3������FΤ���\r_S�J��u1\�<�kX��.>��a��gN�����0B�����u$0��0�}���H./�q�VsD���`qMʛK�X,����K."Xq��TG[�ρ}p-Ձ1=V������_�O���5�[�/kƙ��]���ɋ��{�"Ǉxp;�`h�?�"�Q��ў5\�nE�����ne�����N��UK*�f�7Ӫ�AX���n4r#+Kz�}ձ�%��6v�y���|=�/s���#\� �Y(�xz�����J���0y��o�c@m� >�k���edd�i�R}���@����k��I$Qb
+=�H�͞��u���0 B�7��Eb�[�A���L"��[�]S�8��1��փDQO'~r1��,m�zWw�PoD+���h���*XaY�@'���� �N9m�}W�v����,�J6�J��U�,$j��g�y=�Ϙ-�6���,}X�����S����!3~�Jh���%�5�꟯�!9�2y���$	���
5�Sx��1>[#�ES�f뗇0���]��go��l��ً5��&f�<a�@��
1o�d���fm����[�ݔʣ(���z�.���I3�&fhXlzI�D�#��Y�ے�S�Fps�~�}��������}�j��sܚ�h�p���Gd���*0K�!���h��3~K���<��|j��s�����|]��,h`Ag&u����H-
�	�4Zj������K�5��`���?D?�4	&t85�%�t30Ǯ?q�S����hP�9&�Y��r{�f�`1���� �:R�އPk�\�J�\��#����Ks>�ޘ��9��G�OФb����ԡ���52����Y�jG�c�|�):r&�5{����n:d��G̞$�s�.�s��gR(:���]��^���C7p5��{Q��P�`�S��V�I�I��XA��Y��ns���߮$E�����=�&�s݉պ����,�ʏ
hP�1/WWʍ@��A�,ȡb+����`)������[�{����p�k���Z�T=�+�v�c�f#�)��ֿRޓ	�$_����L$c�����op�-C����iٍ'�ݰ�%��2)6R}�&���;�Y�� �˓�lR����/w&��T~��G>���Fte�>�r&�S���ns����ٔ���OŇ����j�n�H��n& ���x:f��@�$t3�n���F�4SC	gE`�p��T	/w7�����֧�=p�7�$N��FV^�Z��!"��a�
2�j�0T�젅���11���Z|i�3>b�i}���x�v`d��U��%�����������=�O�^_�%ҋ��Г74�r�e�m��~���j��[�8�:Me1BL�J~ר:T���D���J���l�D���#�ki�o[d�y��جSވUmsFc��&�݇k��~R�!��@o�'�h���!+B+\�u��8�3�5bfŶ�11���Ҽ�3�����<`��;SQC��}�1̿��V����d�?g�A�ǰ[�����Bx��N0�,�cp��C�d���
�� �g*I���Pt��5��w���������'p�)uP-�H<	�L#�]��9�_�l�i(��\�'|؃0�2t����l�*"����5�X���Sgf��Ӵ�$l��.T�0iJX�e��W���*^N(�^-#i��^��g3�+j�{��%�vWٳݴ�[z��+#9��Ш]�����Q�Z�J��o��*`���E�?D4�h����Y2 �*=5g݌�)�v,N�cVw�0���HD��2��Ñ����򷄭\甩��7'>Uۀ��G���"7g��^�����SG˚xB%������h��bQ-�)�ֆ��Y�Si��>��,5�>���Ms��s���$�C �1R<0��;q!�������~j����g�d�b*�4n�X���E��T����@U�c���Y�3�ΆJomc���px��g�猥5�]&t#��V}}wZ�2�z�	�q���$M�iq�.��c΋��xw.���'�kM��9�����Î�6G�ؠ�42�{b��Z�s�pu�|O�Lun0�(�޾����ਂ��m�ޫ�Uo7�(v� �W�(s7̈́��v#]ظ9k�T(����|���l$Vm�4����~p�0[���
X��
8���5w��E*bB>AIX(�X��}=?�Ь�~��D��U���w�w!��������F��)т4.&�sy��O���_vR�Y�����5|��0��'w/��r���#� <��N6���|:>��;o����<�z3��wL Y�,��ƕ�S��4ޙ��i�Vk���־UL�J�1��u�U�m�P��3�;h�9�d�r	&�&rN�}�9�h���&᎗�8=tKg@��L��'b��h���'�u��BC���)�����]х�w3��QX�ԧh�ͤʶ�Dv1(VѤϐ��2]�����>W`fy�����3=J��'�g�o5e���*��oHؼ6�N�̮W!�\���d��ɐ�60~7|�s ��#����Ʒ��{{��?��<(C�|bjZq9e��MF�9l��5zn���3q)�I�'AF��{�s�@X뜠Ǥ�KD�r���^���)Ut�ٸ��2�%��=K<I���sM���<3�㣳�H��Ǥ��|x*��5چQ�7�n�4���(�3(!��E��>G7��1��@��h:X��1{ƫ5VV�=��
���W]P�e�Q�C/^Q�g<�ؓ�K���W�HՌJV��¡t$�V����C	�L����x���Ae�:E n�I5�4"���X���p ~¤"H�dk�;7Y��k&������_�Q���%h�+R���Ծ�a穐O���R�?ՉȑN��:����#dr��Ɯ�d"+XV�q'؊��Fx0�!������F����o&��$v�����~Ƃ@���mV;�~�x��w9|#;D>:ןO���^��{��_߉9TcB�����!���#�ͮ��$����7��/������E�����q�dA������cg������+�����6ȕ�Y10a!x�4Hau<.��[�Xs��+7G�$z��/@���&�u�����ynh�D��&�۔����
�!m<W�/ȖīK�uC�K�R (-�߃���f��;����d�Y+���T��X�"L����Y��Nǫ�Z����a� �F�h����s]]*�Ltd�#�J#N��<g��6�(�A�@����N�f�
���X���xx�l랲�_*y>�Ҕ�S���D���I�����V�� �D�J��V+��:Z�>�`�[�����i�d`�k�dlmo���(�� l�~Aln�!��u/��4T\d�G�l���ov!{��U�M���
�`f!�FP�%|o	Рw�3+�F��3y%��F����ƫ4Z3S�p}�Fm�a2#YB�P��͝}t�3#����<��b-�T�ߥ�w��Q.�I+�ru�4����jDw��*&6 �������r7��C"(������fD��E��}�bv�Ic�d�u��&��,j��QޑIO��C(�x�}Q{��@��_g��CF�@��>Ig�#�CJ��63����CU֤՟K3Q���/��ޢ���WL�����	�0�R ���� �L{%��̱5&�0�ҧ��mL$���Ӝ���/ߴ�r��T�u�;{�Q��&T��M��n�>ǖ�Ou5��W��X�Y�*6�N��-��׬�r�!(�!�R�ʍ�u6\2%���ݤ��`	U�N�X��-S�^X�q5��1�f���Cf��OL?����s"9W ��0sC�fU� ��0�B�g����h[n8�b%U��^����i�vb�ԉ�Y�sH�2�[J�+Y��,��x�N/&���,e�YĈ��&�ω�I&�k���-/�RH�2�%RuA��!9���3���,چ����9�)�#Nݐ^IH������Bk�*��u����Zmn}v����r�6�^RɅ ������9��؞ٍH8(R򿈒��,t����-��TaEC�t�� ��E��AЀ9�J�4w����<�@�O�Vah��
���;��֪ngW��Y�p��l�l���S�pB9�qoq}�S�;���{�sMR�<�������W{%_DZ��>� �n��HcK-�?Y��?�L�����x������R�6w�x}���gq��-�/j,���z!/j�S���E���Tg�K�:S�`+�_1�1���V��H�F���3� !�E��>�p�+�̮9�3
��y�?�=k?�`��rpt�T�2�l�~:�BVJ������v��������(���>�o��cp����0q��	�ie�$��F�{�oшx�D��h�B1rʼ��u)�Z�F��83�`�M��Ϋ�ed���kM٥#�4n3 j���}L