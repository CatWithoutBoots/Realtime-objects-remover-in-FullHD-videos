// soc_system_gmm.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module soc_system_gmm (
		input  wire         gmm_fg_detector_cpu_write,      // gmm_fg_detector_cpu.write
		input  wire         gmm_fg_detector_cpu_read,       //                    .read
		input  wire [31:0]  gmm_fg_detector_cpu_writedata,  //                    .writedata
		output wire [31:0]  gmm_fg_detector_cpu_readdata,   //                    .readdata
		input  wire [3:0]   gmm_fg_detector_cpu_address,    //                    .address
		input  wire         gmm_fg_detector_cpu_chipselect, //                    .chipselect
		input  wire [1:0]   gmm_fg_visor_sw_extern,         //     gmm_fg_visor_sw.extern
		input  wire         mem_clk_clk,                    //             mem_clk.clk
		output wire [29:0]  mem_read_address,               //            mem_read.address
		output wire         mem_read_read,                  //                    .read
		output wire [15:0]  mem_read_byteenable,            //                    .byteenable
		input  wire [127:0] mem_read_readdata,              //                    .readdata
		input  wire         mem_read_waitrequest,           //                    .waitrequest
		input  wire         mem_read_readdatavalid,         //                    .readdatavalid
		output wire [6:0]   mem_read_burstcount,            //                    .burstcount
		output wire [29:0]  mem_write_address,              //           mem_write.address
		output wire         mem_write_write,                //                    .write
		output wire [15:0]  mem_write_byteenable,           //                    .byteenable
		output wire [127:0] mem_write_writedata,            //                    .writedata
		input  wire         mem_write_waitrequest,          //                    .waitrequest
		output wire [6:0]   mem_write_burstcount,           //                    .burstcount
		input  wire         rst_reset,                      //                 rst.reset
		input  wire [23:0]  snk_video_data,                 //           snk_video.data
		input  wire         snk_video_endofpacket,          //                    .endofpacket
		output wire         snk_video_ready,                //                    .ready
		input  wire         snk_video_startofpacket,        //                    .startofpacket
		input  wire         snk_video_valid,                //                    .valid
		output wire [23:0]  src_video_data,                 //           src_video.data
		output wire         src_video_endofpacket,          //                    .endofpacket
		input  wire         src_video_ready,                //                    .ready
		output wire         src_video_startofpacket,        //                    .startofpacket
		output wire         src_video_valid                 //                    .valid
	);

	wire   [31:0] gmm_fg_detector_in_pref_readdata;                   // in_dma:prefetcher_csr_readdata -> gmm_fg_detector:in_pref_readdata
	wire    [2:0] gmm_fg_detector_in_pref_address;                    // gmm_fg_detector:in_pref_addr -> in_dma:prefetcher_csr_address
	wire          gmm_fg_detector_in_pref_read;                       // gmm_fg_detector:in_pref_read -> in_dma:prefetcher_csr_read
	wire          gmm_fg_detector_in_pref_write;                      // gmm_fg_detector:in_pref_write -> in_dma:prefetcher_csr_write
	wire   [31:0] gmm_fg_detector_in_pref_writedata;                  // gmm_fg_detector:in_pref_writedata -> in_dma:prefetcher_csr_writedata
	wire   [31:0] gmm_fg_detector_out_pref_readdata;                  // out_dma:prefetcher_csr_readdata -> gmm_fg_detector:out_pref_readdata
	wire    [2:0] gmm_fg_detector_out_pref_address;                   // gmm_fg_detector:out_pref_addr -> out_dma:prefetcher_csr_address
	wire          gmm_fg_detector_out_pref_read;                      // gmm_fg_detector:out_pref_read -> out_dma:prefetcher_csr_read
	wire          gmm_fg_detector_out_pref_write;                     // gmm_fg_detector:out_pref_write -> out_dma:prefetcher_csr_write
	wire   [31:0] gmm_fg_detector_out_pref_writedata;                 // gmm_fg_detector:out_pref_writedata -> out_dma:prefetcher_csr_writedata
	wire          gmm_fg_detector_src_mem_valid;                      // gmm_fg_detector:src_mem_valid -> in_dma:st_sink_valid
	wire  [127:0] gmm_fg_detector_src_mem_data;                       // gmm_fg_detector:src_mem_data -> in_dma:st_sink_data
	wire          gmm_fg_detector_src_mem_ready;                      // in_dma:st_sink_ready -> gmm_fg_detector:src_mem_ready
	wire          gmm_fg_detector_src_mem_startofpacket;              // gmm_fg_detector:src_mem_sop -> in_dma:st_sink_startofpacket
	wire          gmm_fg_detector_src_mem_endofpacket;                // gmm_fg_detector:src_mem_eop -> in_dma:st_sink_endofpacket
	wire    [3:0] gmm_fg_detector_src_mem_empty;                      // gmm_fg_detector:src_mem_empty -> in_dma:st_sink_empty
	wire          gmm_fg_detector_src_video_valid;                    // gmm_fg_detector:src_video_valid -> gmm_fg_visor:snk_valid
	wire   [48:0] gmm_fg_detector_src_video_data;                     // gmm_fg_detector:src_video_data -> gmm_fg_visor:snk_data
	wire          gmm_fg_detector_src_video_ready;                    // gmm_fg_visor:snk_ready -> gmm_fg_detector:src_video_ready
	wire          gmm_fg_detector_src_video_startofpacket;            // gmm_fg_detector:src_video_sop -> gmm_fg_visor:snk_sop
	wire          gmm_fg_detector_src_video_endofpacket;              // gmm_fg_detector:src_video_eop -> gmm_fg_visor:snk_eop
	wire          out_dma_st_source_valid;                            // out_dma:st_source_valid -> gmm_fg_detector:snk_mem_valid
	wire  [127:0] out_dma_st_source_data;                             // out_dma:st_source_data -> gmm_fg_detector:snk_mem_data
	wire          out_dma_st_source_ready;                            // gmm_fg_detector:snk_mem_ready -> out_dma:st_source_ready
	wire          out_dma_st_source_startofpacket;                    // out_dma:st_source_startofpacket -> gmm_fg_detector:snk_mem_sop
	wire          out_dma_st_source_endofpacket;                      // out_dma:st_source_endofpacket -> gmm_fg_detector:snk_mem_eop
	wire    [3:0] out_dma_st_source_empty;                            // out_dma:st_source_empty -> gmm_fg_detector:snk_mem_empty
	wire   [31:0] in_dma_descriptor_read_master_readdata;             // mm_interconnect_0:in_dma_descriptor_read_master_readdata -> in_dma:descriptor_read_master_readdata
	wire          in_dma_descriptor_read_master_waitrequest;          // mm_interconnect_0:in_dma_descriptor_read_master_waitrequest -> in_dma:descriptor_read_master_waitrequest
	wire   [10:0] in_dma_descriptor_read_master_address;              // in_dma:descriptor_read_master_address -> mm_interconnect_0:in_dma_descriptor_read_master_address
	wire          in_dma_descriptor_read_master_read;                 // in_dma:descriptor_read_master_read -> mm_interconnect_0:in_dma_descriptor_read_master_read
	wire          in_dma_descriptor_read_master_readdatavalid;        // mm_interconnect_0:in_dma_descriptor_read_master_readdatavalid -> in_dma:descriptor_read_master_readdatavalid
	wire          in_dma_descriptor_write_master_waitrequest;         // mm_interconnect_0:in_dma_descriptor_write_master_waitrequest -> in_dma:descriptor_write_master_waitrequest
	wire   [10:0] in_dma_descriptor_write_master_address;             // in_dma:descriptor_write_master_address -> mm_interconnect_0:in_dma_descriptor_write_master_address
	wire    [3:0] in_dma_descriptor_write_master_byteenable;          // in_dma:descriptor_write_master_byteenable -> mm_interconnect_0:in_dma_descriptor_write_master_byteenable
	wire    [1:0] in_dma_descriptor_write_master_response;            // mm_interconnect_0:in_dma_descriptor_write_master_response -> in_dma:descriptor_write_master_response
	wire          in_dma_descriptor_write_master_write;               // in_dma:descriptor_write_master_write -> mm_interconnect_0:in_dma_descriptor_write_master_write
	wire   [31:0] in_dma_descriptor_write_master_writedata;           // in_dma:descriptor_write_master_writedata -> mm_interconnect_0:in_dma_descriptor_write_master_writedata
	wire          in_dma_descriptor_write_master_writeresponsevalid;  // mm_interconnect_0:in_dma_descriptor_write_master_writeresponsevalid -> in_dma:descriptor_write_master_writeresponsevalid
	wire          mm_interconnect_0_in_ram_s2_chipselect;             // mm_interconnect_0:in_ram_s2_chipselect -> in_ram:chipselect2
	wire  [255:0] mm_interconnect_0_in_ram_s2_readdata;               // in_ram:readdata2 -> mm_interconnect_0:in_ram_s2_readdata
	wire    [5:0] mm_interconnect_0_in_ram_s2_address;                // mm_interconnect_0:in_ram_s2_address -> in_ram:address2
	wire   [31:0] mm_interconnect_0_in_ram_s2_byteenable;             // mm_interconnect_0:in_ram_s2_byteenable -> in_ram:byteenable2
	wire          mm_interconnect_0_in_ram_s2_write;                  // mm_interconnect_0:in_ram_s2_write -> in_ram:write2
	wire  [255:0] mm_interconnect_0_in_ram_s2_writedata;              // mm_interconnect_0:in_ram_s2_writedata -> in_ram:writedata2
	wire          mm_interconnect_0_in_ram_s2_clken;                  // mm_interconnect_0:in_ram_s2_clken -> in_ram:clken2
	wire   [31:0] out_dma_descriptor_read_master_readdata;            // mm_interconnect_1:out_dma_descriptor_read_master_readdata -> out_dma:descriptor_read_master_readdata
	wire          out_dma_descriptor_read_master_waitrequest;         // mm_interconnect_1:out_dma_descriptor_read_master_waitrequest -> out_dma:descriptor_read_master_waitrequest
	wire   [10:0] out_dma_descriptor_read_master_address;             // out_dma:descriptor_read_master_address -> mm_interconnect_1:out_dma_descriptor_read_master_address
	wire          out_dma_descriptor_read_master_read;                // out_dma:descriptor_read_master_read -> mm_interconnect_1:out_dma_descriptor_read_master_read
	wire          out_dma_descriptor_read_master_readdatavalid;       // mm_interconnect_1:out_dma_descriptor_read_master_readdatavalid -> out_dma:descriptor_read_master_readdatavalid
	wire          out_dma_descriptor_write_master_waitrequest;        // mm_interconnect_1:out_dma_descriptor_write_master_waitrequest -> out_dma:descriptor_write_master_waitrequest
	wire   [10:0] out_dma_descriptor_write_master_address;            // out_dma:descriptor_write_master_address -> mm_interconnect_1:out_dma_descriptor_write_master_address
	wire    [3:0] out_dma_descriptor_write_master_byteenable;         // out_dma:descriptor_write_master_byteenable -> mm_interconnect_1:out_dma_descriptor_write_master_byteenable
	wire    [1:0] out_dma_descriptor_write_master_response;           // mm_interconnect_1:out_dma_descriptor_write_master_response -> out_dma:descriptor_write_master_response
	wire          out_dma_descriptor_write_master_write;              // out_dma:descriptor_write_master_write -> mm_interconnect_1:out_dma_descriptor_write_master_write
	wire   [31:0] out_dma_descriptor_write_master_writedata;          // out_dma:descriptor_write_master_writedata -> mm_interconnect_1:out_dma_descriptor_write_master_writedata
	wire          out_dma_descriptor_write_master_writeresponsevalid; // mm_interconnect_1:out_dma_descriptor_write_master_writeresponsevalid -> out_dma:descriptor_write_master_writeresponsevalid
	wire          mm_interconnect_1_out_ram_s2_chipselect;            // mm_interconnect_1:out_ram_s2_chipselect -> out_ram:chipselect2
	wire  [255:0] mm_interconnect_1_out_ram_s2_readdata;              // out_ram:readdata2 -> mm_interconnect_1:out_ram_s2_readdata
	wire    [5:0] mm_interconnect_1_out_ram_s2_address;               // mm_interconnect_1:out_ram_s2_address -> out_ram:address2
	wire   [31:0] mm_interconnect_1_out_ram_s2_byteenable;            // mm_interconnect_1:out_ram_s2_byteenable -> out_ram:byteenable2
	wire          mm_interconnect_1_out_ram_s2_write;                 // mm_interconnect_1:out_ram_s2_write -> out_ram:write2
	wire  [255:0] mm_interconnect_1_out_ram_s2_writedata;             // mm_interconnect_1:out_ram_s2_writedata -> out_ram:writedata2
	wire          mm_interconnect_1_out_ram_s2_clken;                 // mm_interconnect_1:out_ram_s2_clken -> out_ram:clken2
	wire  [255:0] gmm_fg_detector_in_ram_readdata;                    // mm_interconnect_3:gmm_fg_detector_in_ram_readdata -> gmm_fg_detector:in_ram_readdata
	wire    [5:0] gmm_fg_detector_in_ram_address;                     // gmm_fg_detector:in_ram_addr -> mm_interconnect_3:gmm_fg_detector_in_ram_address
	wire          gmm_fg_detector_in_ram_read;                        // gmm_fg_detector:in_ram_read -> mm_interconnect_3:gmm_fg_detector_in_ram_read
	wire          gmm_fg_detector_in_ram_write;                       // gmm_fg_detector:in_ram_write -> mm_interconnect_3:gmm_fg_detector_in_ram_write
	wire  [255:0] gmm_fg_detector_in_ram_writedata;                   // gmm_fg_detector:in_ram_writedata -> mm_interconnect_3:gmm_fg_detector_in_ram_writedata
	wire          mm_interconnect_3_in_ram_s1_chipselect;             // mm_interconnect_3:in_ram_s1_chipselect -> in_ram:chipselect
	wire  [255:0] mm_interconnect_3_in_ram_s1_readdata;               // in_ram:readdata -> mm_interconnect_3:in_ram_s1_readdata
	wire    [5:0] mm_interconnect_3_in_ram_s1_address;                // mm_interconnect_3:in_ram_s1_address -> in_ram:address
	wire   [31:0] mm_interconnect_3_in_ram_s1_byteenable;             // mm_interconnect_3:in_ram_s1_byteenable -> in_ram:byteenable
	wire          mm_interconnect_3_in_ram_s1_write;                  // mm_interconnect_3:in_ram_s1_write -> in_ram:write
	wire  [255:0] mm_interconnect_3_in_ram_s1_writedata;              // mm_interconnect_3:in_ram_s1_writedata -> in_ram:writedata
	wire          mm_interconnect_3_in_ram_s1_clken;                  // mm_interconnect_3:in_ram_s1_clken -> in_ram:clken
	wire  [255:0] gmm_fg_detector_out_ram_readdata;                   // mm_interconnect_5:gmm_fg_detector_out_ram_readdata -> gmm_fg_detector:out_ram_readdata
	wire    [5:0] gmm_fg_detector_out_ram_address;                    // gmm_fg_detector:out_ram_addr -> mm_interconnect_5:gmm_fg_detector_out_ram_address
	wire          gmm_fg_detector_out_ram_read;                       // gmm_fg_detector:out_ram_read -> mm_interconnect_5:gmm_fg_detector_out_ram_read
	wire          gmm_fg_detector_out_ram_write;                      // gmm_fg_detector:out_ram_write -> mm_interconnect_5:gmm_fg_detector_out_ram_write
	wire  [255:0] gmm_fg_detector_out_ram_writedata;                  // gmm_fg_detector:out_ram_writedata -> mm_interconnect_5:gmm_fg_detector_out_ram_writedata
	wire          mm_interconnect_5_out_ram_s1_chipselect;            // mm_interconnect_5:out_ram_s1_chipselect -> out_ram:chipselect
	wire  [255:0] mm_interconnect_5_out_ram_s1_readdata;              // out_ram:readdata -> mm_interconnect_5:out_ram_s1_readdata
	wire    [5:0] mm_interconnect_5_out_ram_s1_address;               // mm_interconnect_5:out_ram_s1_address -> out_ram:address
	wire   [31:0] mm_interconnect_5_out_ram_s1_byteenable;            // mm_interconnect_5:out_ram_s1_byteenable -> out_ram:byteenable
	wire          mm_interconnect_5_out_ram_s1_write;                 // mm_interconnect_5:out_ram_s1_write -> out_ram:write
	wire  [255:0] mm_interconnect_5_out_ram_s1_writedata;             // mm_interconnect_5:out_ram_s1_writedata -> out_ram:writedata
	wire          mm_interconnect_5_out_ram_s1_clken;                 // mm_interconnect_5:out_ram_s1_clken -> out_ram:clken
	wire          rst_controller_reset_out_reset;                     // rst_controller:reset_out -> [gmm_fg_detector:rst, gmm_fg_visor:rst, in_dma:reset_n_reset_n, in_ram:reset, mm_interconnect_0:in_dma_reset_n_reset_bridge_in_reset_reset, mm_interconnect_1:out_dma_reset_n_reset_bridge_in_reset_reset, mm_interconnect_3:gmm_fg_detector_rst_reset_bridge_in_reset_reset, mm_interconnect_5:gmm_fg_detector_rst_reset_bridge_in_reset_reset, out_dma:reset_n_reset_n, out_ram:reset, rst_translator:in_reset]
	wire          rst_controller_reset_out_reset_req;                 // rst_controller:reset_req -> [in_ram:reset_req, out_ram:reset_req, rst_translator:reset_req_in]

	gmm_fg_detector #(
		.FRAMES_NUM         (2),
		.VIDEO_START_ADDR   (0),
		.VIDEO_SPAN_BYTES   (33177616),
		.CONTROL_SPAN_BYTES (32)
	) gmm_fg_detector (
		.clk                (mem_clk_clk),                             //     clock.clk
		.cpu_write          (gmm_fg_detector_cpu_write),               //       cpu.write
		.cpu_read           (gmm_fg_detector_cpu_read),                //          .read
		.cpu_writedata      (gmm_fg_detector_cpu_writedata),           //          .writedata
		.cpu_readdata       (gmm_fg_detector_cpu_readdata),            //          .readdata
		.cpu_addr           (gmm_fg_detector_cpu_address),             //          .address
		.cpu_cs             (gmm_fg_detector_cpu_chipselect),          //          .chipselect
		.snk_video_data     (snk_video_data),                          // snk_video.data
		.snk_video_eop      (snk_video_endofpacket),                   //          .endofpacket
		.snk_video_ready    (snk_video_ready),                         //          .ready
		.snk_video_sop      (snk_video_startofpacket),                 //          .startofpacket
		.snk_video_valid    (snk_video_valid),                         //          .valid
		.snk_mem_data       (out_dma_st_source_data),                  //   snk_mem.data
		.snk_mem_empty      (out_dma_st_source_empty),                 //          .empty
		.snk_mem_eop        (out_dma_st_source_endofpacket),           //          .endofpacket
		.snk_mem_ready      (out_dma_st_source_ready),                 //          .ready
		.snk_mem_sop        (out_dma_st_source_startofpacket),         //          .startofpacket
		.snk_mem_valid      (out_dma_st_source_valid),                 //          .valid
		.src_video_data     (gmm_fg_detector_src_video_data),          // src_video.data
		.src_video_eop      (gmm_fg_detector_src_video_endofpacket),   //          .endofpacket
		.src_video_ready    (gmm_fg_detector_src_video_ready),         //          .ready
		.src_video_sop      (gmm_fg_detector_src_video_startofpacket), //          .startofpacket
		.src_video_valid    (gmm_fg_detector_src_video_valid),         //          .valid
		.src_mem_data       (gmm_fg_detector_src_mem_data),            //   src_mem.data
		.src_mem_empty      (gmm_fg_detector_src_mem_empty),           //          .empty
		.src_mem_eop        (gmm_fg_detector_src_mem_endofpacket),     //          .endofpacket
		.src_mem_ready      (gmm_fg_detector_src_mem_ready),           //          .ready
		.src_mem_sop        (gmm_fg_detector_src_mem_startofpacket),   //          .startofpacket
		.src_mem_valid      (gmm_fg_detector_src_mem_valid),           //          .valid
		.rst                (rst_controller_reset_out_reset),          //       rst.reset
		.in_ram_addr        (gmm_fg_detector_in_ram_address),          //    in_ram.address
		.in_ram_write       (gmm_fg_detector_in_ram_write),            //          .write
		.in_ram_writedata   (gmm_fg_detector_in_ram_writedata),        //          .writedata
		.in_ram_read        (gmm_fg_detector_in_ram_read),             //          .read
		.in_ram_readdata    (gmm_fg_detector_in_ram_readdata),         //          .readdata
		.out_ram_addr       (gmm_fg_detector_out_ram_address),         //   out_ram.address
		.out_ram_write      (gmm_fg_detector_out_ram_write),           //          .write
		.out_ram_writedata  (gmm_fg_detector_out_ram_writedata),       //          .writedata
		.out_ram_read       (gmm_fg_detector_out_ram_read),            //          .read
		.out_ram_readdata   (gmm_fg_detector_out_ram_readdata),        //          .readdata
		.in_pref_addr       (gmm_fg_detector_in_pref_address),         //   in_pref.address
		.in_pref_write      (gmm_fg_detector_in_pref_write),           //          .write
		.in_pref_writedata  (gmm_fg_detector_in_pref_writedata),       //          .writedata
		.in_pref_read       (gmm_fg_detector_in_pref_read),            //          .read
		.in_pref_readdata   (gmm_fg_detector_in_pref_readdata),        //          .readdata
		.out_pref_addr      (gmm_fg_detector_out_pref_address),        //  out_pref.address
		.out_pref_write     (gmm_fg_detector_out_pref_write),          //          .write
		.out_pref_writedata (gmm_fg_detector_out_pref_writedata),      //          .writedata
		.out_pref_read      (gmm_fg_detector_out_pref_read),           //          .read
		.out_pref_readdata  (gmm_fg_detector_out_pref_readdata)        //          .readdata
	);

	gmm_fg_visor gmm_fg_visor (
		.rst       (rst_controller_reset_out_reset),          // rst.reset
		.clk       (mem_clk_clk),                             // clk.clk
		.snk_data  (gmm_fg_detector_src_video_data),          // snk.data
		.snk_eop   (gmm_fg_detector_src_video_endofpacket),   //    .endofpacket
		.snk_ready (gmm_fg_detector_src_video_ready),         //    .ready
		.snk_sop   (gmm_fg_detector_src_video_startofpacket), //    .startofpacket
		.snk_valid (gmm_fg_detector_src_video_valid),         //    .valid
		.src_data  (src_video_data),                          // src.data
		.src_eop   (src_video_endofpacket),                   //    .endofpacket
		.src_ready (src_video_ready),                         //    .ready
		.src_sop   (src_video_startofpacket),                 //    .startofpacket
		.src_valid (src_video_valid),                         //    .valid
		.sw        (gmm_fg_visor_sw_extern)                   //  sw.extern
	);

	soc_system_gmm_in_dma in_dma (
		.mm_write_address                           (mem_write_address),                                 //                mm_write.address
		.mm_write_write                             (mem_write_write),                                   //                        .write
		.mm_write_byteenable                        (mem_write_byteenable),                              //                        .byteenable
		.mm_write_writedata                         (mem_write_writedata),                               //                        .writedata
		.mm_write_waitrequest                       (mem_write_waitrequest),                             //                        .waitrequest
		.mm_write_burstcount                        (mem_write_burstcount),                              //                        .burstcount
		.descriptor_read_master_address             (in_dma_descriptor_read_master_address),             //  descriptor_read_master.address
		.descriptor_read_master_read                (in_dma_descriptor_read_master_read),                //                        .read
		.descriptor_read_master_readdata            (in_dma_descriptor_read_master_readdata),            //                        .readdata
		.descriptor_read_master_waitrequest         (in_dma_descriptor_read_master_waitrequest),         //                        .waitrequest
		.descriptor_read_master_readdatavalid       (in_dma_descriptor_read_master_readdatavalid),       //                        .readdatavalid
		.descriptor_write_master_address            (in_dma_descriptor_write_master_address),            // descriptor_write_master.address
		.descriptor_write_master_write              (in_dma_descriptor_write_master_write),              //                        .write
		.descriptor_write_master_byteenable         (in_dma_descriptor_write_master_byteenable),         //                        .byteenable
		.descriptor_write_master_writedata          (in_dma_descriptor_write_master_writedata),          //                        .writedata
		.descriptor_write_master_waitrequest        (in_dma_descriptor_write_master_waitrequest),        //                        .waitrequest
		.descriptor_write_master_response           (in_dma_descriptor_write_master_response),           //                        .response
		.descriptor_write_master_writeresponsevalid (in_dma_descriptor_write_master_writeresponsevalid), //                        .writeresponsevalid
		.clock_clk                                  (mem_clk_clk),                                       //                   clock.clk
		.reset_n_reset_n                            (~rst_controller_reset_out_reset),                   //                 reset_n.reset_n
		.csr_writedata                              (),                                                  //                     csr.writedata
		.csr_write                                  (),                                                  //                        .write
		.csr_byteenable                             (),                                                  //                        .byteenable
		.csr_readdata                               (),                                                  //                        .readdata
		.csr_read                                   (),                                                  //                        .read
		.csr_address                                (),                                                  //                        .address
		.prefetcher_csr_address                     (gmm_fg_detector_in_pref_address),                   //          prefetcher_csr.address
		.prefetcher_csr_read                        (gmm_fg_detector_in_pref_read),                      //                        .read
		.prefetcher_csr_write                       (gmm_fg_detector_in_pref_write),                     //                        .write
		.prefetcher_csr_writedata                   (gmm_fg_detector_in_pref_writedata),                 //                        .writedata
		.prefetcher_csr_readdata                    (gmm_fg_detector_in_pref_readdata),                  //                        .readdata
		.csr_irq_irq                                (),                                                  //                 csr_irq.irq
		.st_sink_data                               (gmm_fg_detector_src_mem_data),                      //                 st_sink.data
		.st_sink_valid                              (gmm_fg_detector_src_mem_valid),                     //                        .valid
		.st_sink_ready                              (gmm_fg_detector_src_mem_ready),                     //                        .ready
		.st_sink_startofpacket                      (gmm_fg_detector_src_mem_startofpacket),             //                        .startofpacket
		.st_sink_endofpacket                        (gmm_fg_detector_src_mem_endofpacket),               //                        .endofpacket
		.st_sink_empty                              (gmm_fg_detector_src_mem_empty)                      //                        .empty
	);

	soc_system_gmm_in_ram in_ram (
		.address     (mm_interconnect_3_in_ram_s1_address),    //     s1.address
		.clken       (mm_interconnect_3_in_ram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_3_in_ram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_3_in_ram_s1_write),      //       .write
		.readdata    (mm_interconnect_3_in_ram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_3_in_ram_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_3_in_ram_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_0_in_ram_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_in_ram_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_in_ram_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_in_ram_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_in_ram_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_in_ram_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_in_ram_s2_byteenable), //       .byteenable
		.clk         (mem_clk_clk),                            //   clk1.clk
		.reset       (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),     //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	soc_system_gmm_out_dma out_dma (
		.mm_read_address                            (mem_read_address),                                   //                 mm_read.address
		.mm_read_read                               (mem_read_read),                                      //                        .read
		.mm_read_byteenable                         (mem_read_byteenable),                                //                        .byteenable
		.mm_read_readdata                           (mem_read_readdata),                                  //                        .readdata
		.mm_read_waitrequest                        (mem_read_waitrequest),                               //                        .waitrequest
		.mm_read_readdatavalid                      (mem_read_readdatavalid),                             //                        .readdatavalid
		.mm_read_burstcount                         (mem_read_burstcount),                                //                        .burstcount
		.descriptor_read_master_address             (out_dma_descriptor_read_master_address),             //  descriptor_read_master.address
		.descriptor_read_master_read                (out_dma_descriptor_read_master_read),                //                        .read
		.descriptor_read_master_readdata            (out_dma_descriptor_read_master_readdata),            //                        .readdata
		.descriptor_read_master_waitrequest         (out_dma_descriptor_read_master_waitrequest),         //                        .waitrequest
		.descriptor_read_master_readdatavalid       (out_dma_descriptor_read_master_readdatavalid),       //                        .readdatavalid
		.descriptor_write_master_address            (out_dma_descriptor_write_master_address),            // descriptor_write_master.address
		.descriptor_write_master_write              (out_dma_descriptor_write_master_write),              //                        .write
		.descriptor_write_master_byteenable         (out_dma_descriptor_write_master_byteenable),         //                        .byteenable
		.descriptor_write_master_writedata          (out_dma_descriptor_write_master_writedata),          //                        .writedata
		.descriptor_write_master_waitrequest        (out_dma_descriptor_write_master_waitrequest),        //                        .waitrequest
		.descriptor_write_master_response           (out_dma_descriptor_write_master_response),           //                        .response
		.descriptor_write_master_writeresponsevalid (out_dma_descriptor_write_master_writeresponsevalid), //                        .writeresponsevalid
		.clock_clk                                  (mem_clk_clk),                                        //                   clock.clk
		.reset_n_reset_n                            (~rst_controller_reset_out_reset),                    //                 reset_n.reset_n
		.csr_writedata                              (),                                                   //                     csr.writedata
		.csr_write                                  (),                                                   //                        .write
		.csr_byteenable                             (),                                                   //                        .byteenable
		.csr_readdata                               (),                                                   //                        .readdata
		.csr_read                                   (),                                                   //                        .read
		.csr_address                                (),                                                   //                        .address
		.prefetcher_csr_address                     (gmm_fg_detector_out_pref_address),                   //          prefetcher_csr.address
		.prefetcher_csr_read                        (gmm_fg_detector_out_pref_read),                      //                        .read
		.prefetcher_csr_write                       (gmm_fg_detector_out_pref_write),                     //                        .write
		.prefetcher_csr_writedata                   (gmm_fg_detector_out_pref_writedata),                 //                        .writedata
		.prefetcher_csr_readdata                    (gmm_fg_detector_out_pref_readdata),                  //                        .readdata
		.csr_irq_irq                                (),                                                   //                 csr_irq.irq
		.st_source_data                             (out_dma_st_source_data),                             //               st_source.data
		.st_source_valid                            (out_dma_st_source_valid),                            //                        .valid
		.st_source_ready                            (out_dma_st_source_ready),                            //                        .ready
		.st_source_startofpacket                    (out_dma_st_source_startofpacket),                    //                        .startofpacket
		.st_source_endofpacket                      (out_dma_st_source_endofpacket),                      //                        .endofpacket
		.st_source_empty                            (out_dma_st_source_empty)                             //                        .empty
	);

	soc_system_gmm_out_ram out_ram (
		.address     (mm_interconnect_5_out_ram_s1_address),    //     s1.address
		.clken       (mm_interconnect_5_out_ram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_5_out_ram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_5_out_ram_s1_write),      //       .write
		.readdata    (mm_interconnect_5_out_ram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_5_out_ram_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_5_out_ram_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_1_out_ram_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_1_out_ram_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_1_out_ram_s2_clken),      //       .clken
		.write2      (mm_interconnect_1_out_ram_s2_write),      //       .write
		.readdata2   (mm_interconnect_1_out_ram_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_1_out_ram_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_1_out_ram_s2_byteenable), //       .byteenable
		.clk         (mem_clk_clk),                             //   clk1.clk
		.reset       (rst_controller_reset_out_reset),          // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),      //       .reset_req
		.freeze      (1'b0)                                     // (terminated)
	);

	soc_system_gmm_mm_interconnect_0 mm_interconnect_0 (
		.mem_clk_out_clk_clk                               (mem_clk_clk),                                       //                      mem_clk_out_clk.clk
		.in_dma_reset_n_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                    // in_dma_reset_n_reset_bridge_in_reset.reset
		.in_dma_descriptor_read_master_address             (in_dma_descriptor_read_master_address),             //        in_dma_descriptor_read_master.address
		.in_dma_descriptor_read_master_waitrequest         (in_dma_descriptor_read_master_waitrequest),         //                                     .waitrequest
		.in_dma_descriptor_read_master_read                (in_dma_descriptor_read_master_read),                //                                     .read
		.in_dma_descriptor_read_master_readdata            (in_dma_descriptor_read_master_readdata),            //                                     .readdata
		.in_dma_descriptor_read_master_readdatavalid       (in_dma_descriptor_read_master_readdatavalid),       //                                     .readdatavalid
		.in_dma_descriptor_write_master_address            (in_dma_descriptor_write_master_address),            //       in_dma_descriptor_write_master.address
		.in_dma_descriptor_write_master_waitrequest        (in_dma_descriptor_write_master_waitrequest),        //                                     .waitrequest
		.in_dma_descriptor_write_master_byteenable         (in_dma_descriptor_write_master_byteenable),         //                                     .byteenable
		.in_dma_descriptor_write_master_write              (in_dma_descriptor_write_master_write),              //                                     .write
		.in_dma_descriptor_write_master_writedata          (in_dma_descriptor_write_master_writedata),          //                                     .writedata
		.in_dma_descriptor_write_master_response           (in_dma_descriptor_write_master_response),           //                                     .response
		.in_dma_descriptor_write_master_writeresponsevalid (in_dma_descriptor_write_master_writeresponsevalid), //                                     .writeresponsevalid
		.in_ram_s2_address                                 (mm_interconnect_0_in_ram_s2_address),               //                            in_ram_s2.address
		.in_ram_s2_write                                   (mm_interconnect_0_in_ram_s2_write),                 //                                     .write
		.in_ram_s2_readdata                                (mm_interconnect_0_in_ram_s2_readdata),              //                                     .readdata
		.in_ram_s2_writedata                               (mm_interconnect_0_in_ram_s2_writedata),             //                                     .writedata
		.in_ram_s2_byteenable                              (mm_interconnect_0_in_ram_s2_byteenable),            //                                     .byteenable
		.in_ram_s2_chipselect                              (mm_interconnect_0_in_ram_s2_chipselect),            //                                     .chipselect
		.in_ram_s2_clken                                   (mm_interconnect_0_in_ram_s2_clken)                  //                                     .clken
	);

	soc_system_gmm_mm_interconnect_1 mm_interconnect_1 (
		.mem_clk_out_clk_clk                                (mem_clk_clk),                                        //                       mem_clk_out_clk.clk
		.out_dma_reset_n_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                     // out_dma_reset_n_reset_bridge_in_reset.reset
		.out_dma_descriptor_read_master_address             (out_dma_descriptor_read_master_address),             //        out_dma_descriptor_read_master.address
		.out_dma_descriptor_read_master_waitrequest         (out_dma_descriptor_read_master_waitrequest),         //                                      .waitrequest
		.out_dma_descriptor_read_master_read                (out_dma_descriptor_read_master_read),                //                                      .read
		.out_dma_descriptor_read_master_readdata            (out_dma_descriptor_read_master_readdata),            //                                      .readdata
		.out_dma_descriptor_read_master_readdatavalid       (out_dma_descriptor_read_master_readdatavalid),       //                                      .readdatavalid
		.out_dma_descriptor_write_master_address            (out_dma_descriptor_write_master_address),            //       out_dma_descriptor_write_master.address
		.out_dma_descriptor_write_master_waitrequest        (out_dma_descriptor_write_master_waitrequest),        //                                      .waitrequest
		.out_dma_descriptor_write_master_byteenable         (out_dma_descriptor_write_master_byteenable),         //                                      .byteenable
		.out_dma_descriptor_write_master_write              (out_dma_descriptor_write_master_write),              //                                      .write
		.out_dma_descriptor_write_master_writedata          (out_dma_descriptor_write_master_writedata),          //                                      .writedata
		.out_dma_descriptor_write_master_response           (out_dma_descriptor_write_master_response),           //                                      .response
		.out_dma_descriptor_write_master_writeresponsevalid (out_dma_descriptor_write_master_writeresponsevalid), //                                      .writeresponsevalid
		.out_ram_s2_address                                 (mm_interconnect_1_out_ram_s2_address),               //                            out_ram_s2.address
		.out_ram_s2_write                                   (mm_interconnect_1_out_ram_s2_write),                 //                                      .write
		.out_ram_s2_readdata                                (mm_interconnect_1_out_ram_s2_readdata),              //                                      .readdata
		.out_ram_s2_writedata                               (mm_interconnect_1_out_ram_s2_writedata),             //                                      .writedata
		.out_ram_s2_byteenable                              (mm_interconnect_1_out_ram_s2_byteenable),            //                                      .byteenable
		.out_ram_s2_chipselect                              (mm_interconnect_1_out_ram_s2_chipselect),            //                                      .chipselect
		.out_ram_s2_clken                                   (mm_interconnect_1_out_ram_s2_clken)                  //                                      .clken
	);

	soc_system_gmm_mm_interconnect_3 mm_interconnect_3 (
		.mem_clk_out_clk_clk                             (mem_clk_clk),                            //                           mem_clk_out_clk.clk
		.gmm_fg_detector_rst_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),         // gmm_fg_detector_rst_reset_bridge_in_reset.reset
		.gmm_fg_detector_in_ram_address                  (gmm_fg_detector_in_ram_address),         //                    gmm_fg_detector_in_ram.address
		.gmm_fg_detector_in_ram_read                     (gmm_fg_detector_in_ram_read),            //                                          .read
		.gmm_fg_detector_in_ram_readdata                 (gmm_fg_detector_in_ram_readdata),        //                                          .readdata
		.gmm_fg_detector_in_ram_write                    (gmm_fg_detector_in_ram_write),           //                                          .write
		.gmm_fg_detector_in_ram_writedata                (gmm_fg_detector_in_ram_writedata),       //                                          .writedata
		.in_ram_s1_address                               (mm_interconnect_3_in_ram_s1_address),    //                                 in_ram_s1.address
		.in_ram_s1_write                                 (mm_interconnect_3_in_ram_s1_write),      //                                          .write
		.in_ram_s1_readdata                              (mm_interconnect_3_in_ram_s1_readdata),   //                                          .readdata
		.in_ram_s1_writedata                             (mm_interconnect_3_in_ram_s1_writedata),  //                                          .writedata
		.in_ram_s1_byteenable                            (mm_interconnect_3_in_ram_s1_byteenable), //                                          .byteenable
		.in_ram_s1_chipselect                            (mm_interconnect_3_in_ram_s1_chipselect), //                                          .chipselect
		.in_ram_s1_clken                                 (mm_interconnect_3_in_ram_s1_clken)       //                                          .clken
	);

	soc_system_gmm_mm_interconnect_5 mm_interconnect_5 (
		.mem_clk_out_clk_clk                             (mem_clk_clk),                             //                           mem_clk_out_clk.clk
		.gmm_fg_detector_rst_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),          // gmm_fg_detector_rst_reset_bridge_in_reset.reset
		.gmm_fg_detector_out_ram_address                 (gmm_fg_detector_out_ram_address),         //                   gmm_fg_detector_out_ram.address
		.gmm_fg_detector_out_ram_read                    (gmm_fg_detector_out_ram_read),            //                                          .read
		.gmm_fg_detector_out_ram_readdata                (gmm_fg_detector_out_ram_readdata),        //                                          .readdata
		.gmm_fg_detector_out_ram_write                   (gmm_fg_detector_out_ram_write),           //                                          .write
		.gmm_fg_detector_out_ram_writedata               (gmm_fg_detector_out_ram_writedata),       //                                          .writedata
		.out_ram_s1_address                              (mm_interconnect_5_out_ram_s1_address),    //                                out_ram_s1.address
		.out_ram_s1_write                                (mm_interconnect_5_out_ram_s1_write),      //                                          .write
		.out_ram_s1_readdata                             (mm_interconnect_5_out_ram_s1_readdata),   //                                          .readdata
		.out_ram_s1_writedata                            (mm_interconnect_5_out_ram_s1_writedata),  //                                          .writedata
		.out_ram_s1_byteenable                           (mm_interconnect_5_out_ram_s1_byteenable), //                                          .byteenable
		.out_ram_s1_chipselect                           (mm_interconnect_5_out_ram_s1_chipselect), //                                          .chipselect
		.out_ram_s1_clken                                (mm_interconnect_5_out_ram_s1_clken)       //                                          .clken
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (rst_reset),                          // reset_in0.reset
		.clk            (mem_clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
