��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&��^L�h�m��uXҰ��>�!Ə�)V?9�d@:	P�Y���������٫�(59Au[�n�!.I1?�Ĭ�<��6&+:���7�I��!���!��~cq����8B��-ս��P��P�z�M-�@7X�ˏ[�OX�"�,��m� ;e��u��W[�J�A�G�G��"GU�7��%�a���F�{zV�4ː��A�WX9�4,��P��G�-��\o�#U�{Rמjr��as0�a����#~�b_��D&=��]�V׆(ͩ�eh.(c�XT�s`l��P�+c��bS|��폐��L�\�n?�8��f��r�3���x�Q�ZZA\se�e�9ViL4:XA7�k4�~3Y~�FS~��w�U�!�eX���Cj��H���DѤ���b⾮�~걚�I�3��<j.1�b�!����y�ӣ���<'�k��Yҁ�`g2���0�Z�{��j��j����g���!��C[�,���<������'�o�� r)�FH�c�ץ�s��T��B�Fg
�I�J�9hw�F���z�5M��ݰ�h�=�K�J�f��sr������Y;��=�iM���hV(�=�|_�`������
X8�b�+Z�	��c0=N�E�R�ɖ2�pTn�fP5��y+��b�����1>)��2��jD� z�f]��&=Մ�@������V�U.�e .M~���Kj��G����_Є�S������6�w��A���r�����QЧև6���w��uL.�nP�Ж
��w�8��s�A���~��#�䧁���
���Ѽ8�	(x�c��q)��&a\}�~+��9�3]���'�����?\Ys���~��7c{�y��7�Wڼ@g�`Mz��D���w���3��{��?�ְ�
�D]��@���5
������R����_Ī��8�&W}�xȬ&c	����X�EZd����g�2�9W|6�&�a�����C9;�7(3�ڵr-ݴ�5��?�̃�Cm��D��0�e~q����x���z�ڟH?�]��e9��>� �����k}���U���j;��;���h����Ŝ$�aؒ8r^ �y�Z�օGƃP�1�O'8�(��_ f������iG�tLf���@��D��(�r�;��Qk�[�KvR6��\�tK%���2���w�9ib�F��w�2���9�_���m�^�-*����R�[<9U\�U���4ʵjK�	�J&�m!s����x�W�����u�\9 24�vʑĄt���)v�#.�`����q ���?f�v!���eBA���ۻ ᵗ�F�A�s\	�����FI٘����*	��٭�p_:t	���h�}�oC2.�ws�8�Y�3���N�T��ʘ�f���Ҩµo)��=5@�T-gc��M�xg����[l'.����y{cF��9��]�����6K
�J��EC�Zڝi���:kH����:0��E�y}0�n����)�6�Ҭ�q��Y:��vٯ���k7K]q 6D�)�Hi�����x��?q����6�w^�Y��Tl�w� "��AL;7OM����W~�M���P���O�͟�������tȃk�|�0J��k4?H"p���7��8[��&H�k�}�e���F2�_ߺ��2[4��Y	��m�'�镘��'��C��P�d�ҳ���i�ZnZ���?�o"��~6ʱajȒ���1?rR2�u7Ӝ�H����|�Ǽj/��+�ӻ���	H����@���?�c{���������H89@���>�)N1��1%R�s���-%��K>e3��O���:h7r)��+1�O7zR#���O�nQ��

�(r��:�Qb*$=��?�����gmm�sJ��`�k��ązG�0�Ӳ�؋�˄�Pw����U[�P���2�U2"3��y�2.KK}����¡}=�媺U��h�_� ���uX<��ۗ��'r�*���v���C���z��!jvщ��TP��Y���,ܩT8BT�._���9
�䒚��%v`8H�>����,�i}�<I���B�"T��t�����w(:ޜE s�M��o	6;j'�����+v�L�J$��~�$�U(s'��C�Ѱ樖�[�_��_V��"b���s�x7o��?�sp,:�Q:	�D߉y\��_��k&�ȳ|�w�s����i� ��7�������VX��WR��^e��8.oHw�|2K��:���P5�E���Y>��u%�d��'駇���X���la[�y�{�K�r�2��)p�*?�����:92{�`:���S�z2�"B�vލ'NE��R!u�XT�:ݮ��$�Rx���vV�� ��ۃVz�'�{e	�gi�c0m�Q��+1[�u~��Sǻ�_�=8���=	j��j�u��L�~i�
�e����Q��ٖ0*+�v(�h1���
V����~SBƶ�������L����1�������,��!��5k�Nw��U'q�X'���D."d���J���Q����9���s$J'��6�C�a�-!*8��gj���%m���SNY�4U�ϭ��V]\��|�B��-��[��Dq�O�ɐ�KVx5EYn W8����-�C�׻��_���Ff:�����ܦ2,��[)�g'�2�!�(�X�?�	k�g��֌Ur3�Z���
�3�����с��|��+P�` ��mG�rG��gO�IX����*?��=�c�x���(������΋{���'ݮ����؀��%�Y����)�Ώ�[С?���k�|$+9��t����O�W�m(�{"S���&!T<��	�11hzGIf��ˍ�j!���;	�͡��f:^�:P��x�Oi<��2A�aA�X�Fv�����uT���ɱ�s{��D�(���ZRZE�I�jƍ�8<�1rn+�����M�I9��:�
W����lQ�!6n��z�)|����#�Յo�0n@v꧁p.	d!�tq%-�<�)���y~M~-�tY�^���&"�X��Y{􃳻��$E_�WI`���`C;
L�
�l��k�;�ϭ�}��-+���F*���*����?�`��0��Ҋ(��z�ep��Kx'vY�^/���_�yI�08�3W
(��[�&Ӟ�4k^S��c�9��N��ǎ�.�y��l*��Z)�_�����<hС�ڙ@���>��MP���G������H�1jD�
Cx@4��@�	HԠ�P}YPC��q�:rj���_��S�$>�8D��6������^�
Ȃ��, �u��i6LW�̴��hӃ֞S��6����Xwc�K�M����z�l�.�缩�7z-��	����7ԹB�̫#�,�[��	5h�=Zܬ
�
X�pi��)��3X��:��CD�t�M�v�����D�`�(�GS�i��]n*jCݟs���?a~�y���P��ӕ5-�s�G?#��8�yIA����@��4���ur\Y|�Xe+�RBN�� U��,Z��i���oB/2�z�3F��7L$��9H��Y��/��U3
�?%sV=��P�N�@1O62��b�Q��!|�A�&�E]T){�m� ��*?�E��G+>s�Z�n�i�t�X1v�uRr��Ķu(�S.s�L3�Rt���Mՠ�
� �1���.v�@ٴTS��#��z*1�2�H3<�z$�~v��Lv'�\�����:7MH�^/���?�������;&�Du��X�u&��[�����l`D,�f� @���n�;���÷�f�;&\NIu�� ��1�;��Ҙ*5�|@���L��0`�j�� �eωeb�M��R)��i�hfv��8p�Z:L�{;f� �ʀѽ�K�y /3�E�Y�.�b�!���� a{M��q�Q<K�r<w� @�D�
�U�xEhQ���?%K�!Y�گ�[�_�W�v�`b��,J4�
L*�<�+��#���Z����D4�n�@J��&x�i�f��d5XFK�G�����)�S�EË�?8��3�J YV�Z�<	}��XϩyZ@��c-�ϥ�+ʍ�p����a�stSb�ઘ�+�l8߄����=[)峇���~u؝��d����b�E\���}b�9��2�W@��[������x�؉2r-�}��t��i5�s��s�z�>���o�8��a{ԝ��Y�+�@$P�a��]�� K�y"��A���	����j�%�:\P��c��V�4�8ƌ�<��`{^nP����\$ή/�O>�sμ�Ⱦ6ῶo�#��x�^J,��va��I뚱e����[�n�|I|�/�q\Ԡ�Y�t1��ߎ�s�|_s�c~��;�H�����2��^�*�V��B�ύ�i���r�T�WL��s
����e�\�N߿�&b��m�6��`�h��M^c���r3��3�����k����ߤo ������bRQl�;��s�	�w�|$�喙h%�8f.���Y���F����7����&�nb997S�ƎNw���8e>�>؄��;��d�j:b�ߗC��Aw]�It�~)�EEO'O��O��SP�����AN���£&!��.���� 0�=� �F�"Ø�j��(�fI=�nx��+1�=e#���U=}dV�1&J�Tu�oG���x��R����,�m��{�YJ��m�N�x�Ss?�������mc�zm�w@��!R��ؾ_�*a�������xq��^��$���\�Z�v�F��Bد�4���6����t�t?�҈�F�;PiU�8;Q=.0E��'��e�,v�����y��J�N�����5^i�l��\Г%g���7$5���l�ڻ!-�<t��̤rU�mZ��ΝM�?LZ���O����e�C��{�i��|��v �������<w���9���̇V����4�3��I�~q�R��|�ֻnM�o�������~CE~E���S�w�q�Ʉ}��I��!��bVm�޾P�ED����e}յ���س�I��U�5�o��y4��aqbxW����e���k� ��:�II^{&���qa~Y("1-�I���uR�̣ J*�e����F������[_%h�?���\�:3��s��OV�)_�I�^_�9��99�����Z�(�K�PF��=,+�K]�"�䕝I�������� :�����{�+>����s��6�3�>d�� Y���;Xr����d��J6T=�X�^�6��4L{^��[�6u����!��1�g��N-,k�]�-�+
B�=|��\_0(�1�0	��9�6R\���L"�����4��ȫb{&1�VW?-���S�{KK���'WQ"L�+7��( �(K.f��Si��EΤ �i�+)�K��� ^�Ά�J�����>|���,bu�@�?~��I�ڲ���C�e�Շ���Vk�?{0�܇w���g�(�ոkė��B�/�ɕ�ܼF�SW�9�*S:� �i6ZN�9�����x�e*�]�U�k!$��0UԦЊ������(gעX�1n��g�Xy�m��xy�@��B>;�e.��~m���Y�Aj���y�~��0#�W���Mf���B�+��]C�c7cBF3<��&v��"6&gV u)��SKg_:�(�� �U�`7��r
.K��pyG�2�fo��r;X��62B��@��K� ������Β@�y��]��j�e�����kg��J�4O��42��X�;P�d�W�-%+&��E��߄0��rmc���vpzY�8�d��EH�Y�F�	I��ݒHҝ�SC��e�1�#$@�q���<E��� Ԇ;��N�W�n����ꊋE\Kmk����0}�6��BY�.��#E��13�� O5��pt#�|�Og�74�
�J��4�`��E͋��	�P,F稛��o/䶧%|O�PC8����? 1����q+V�wC�J6��&��a�V��Ý�Su�1oovfO7MV~��Z�,�a8��&q�c�?T�O�8�`��}c�P�,�Fy����^C�
,�(:'���sa����ф����Ȭ��^�-n�ȊT�P�e���2�7�F����+����H��Ӱ�#ﱩ�'����#��/��f�]����\�Mϔ/��P�n8���w�-�@y�I��y�#����v_b��sy��|ڨ��/QIA*�|��� �Y���9|r�T�ӹ�緩�1�y]��A||�`�C������ vc�6ι�.J[�U֖G6	F�P��oam�ȱZ�"���	���#�x�X��C�6;f�ՃQƶ�2$}_�A�Hk���~GP9 _��=��M�B��@���g�ǶK "=�eO�����1g��������V]�߲�g,�i�Dy1v
+�s� �S�C���B8�pc^ɪ�H�ג�	!�y�[�T	�b`u�mh�uL+tO�Z��8Ӆ1�4T5�\8*�V2{#X�����R�CZέ�.՞��՚Ҷ�r",�ȑ7}�� ���c}�v6\����q[[P<��J1.�sȤTH���ǮKK
Vt�OH�7	�j�Y�ʺ��C����+r�xv��E�*�� #������"�1&mʳ�Y�q���9���Z�o��:��"Vɛ�K�]��x�,�[��Nl�:D+Z�\��P�������*���Uvih��ll��P�
*�	�V(�aF2V������[^���T�;���Wc*clh�,Bi��g�Zr_?Lx��k?�:Hl"�P#0PY���,�~�w	r��5hc��](uG��T �yYS��*���������0̖��ڌ��z��d9�>���-��uY���hLٲٝʹ���Р�\\�{�n��2��B��p�
����,�%9( �-~�t�,#(�"��i�F���`n��-5^�)��ƫB�"��}Zz��i���r��&±|��(�M����2G<ctXk(��JGG�:��N�d'�JlV�y����I���#@�W\��:Gr\��&�������e"���l�
ɇ��>v �G�n
-a�kDNXm��I���Yl�mXds�Ђ�7y�.V(��E?�<W�1O��񏃹;�h�p9�n�S|�`q���TʙD1��?D�H�Ē����E�g�i1��-��׾V���]�/"3ҝ��ζ�����-����ak?bba�A;HZ�B�9-�<ɠ,�n5~�Y��30(О2�y�?�ѷg��J�C�0ؾ,o��GQK��>{JM�j����X���?*2�� ��E_b(
��_)�O�/'H���R��)�E^��@x��YT���$�� h��V��܌��D��Ē�?T>���g�S�	�gtNDկtѸ��
�*�oR��"�,+n�6f��x)�B9,���@V�A��+w�Y�p"qs�!�,h���yV�B��� &��ׁzkjM>�[�C��d����""kVd"��J�K�1���WlQ�f��-<�I
��I	���*�٥�>����Y�W�R6p�%*���q<cEt<Z
��`����Stz�cQ3y��D-ǅj:���6���$�Ե�
����X�=e4`� �Fb�3N��#͑2��W�	�Zʔ:]�eh�V#��Cu.�v���?�y29�xm�a�Ε�m����PRZ{�h"�<Cz	�8���L��]
�kV%%*J{z:���_U��R��!�$�������4�ݢ�w8ҋ|��.��"�*�]k���p��������A�>O ��.|�pN9U�\����t�2g߾g/���bJ�����75)r�=H)����ChM��jd��p=c��� �9�A��"G�Z�[b�meb�K�����8
}��m׽�M�MY���ެ�(���9X|>�� �Ib4�I@�|`���Z�:���� _:�r��'7����)"�_��U�_H��[EB|�2ONq���#��������K�0�rX>�M8��@�"G�2&ٞ"(�=�tC$P��O� u_ ��~�L�B��8�a�/�}nI�&�hL�7��m�h��9���ϵ�>۰|�$��)��6r~�of@~�b*GӢG0z8�S�����[�W�[���)��F�#%QC�� =g�O�4/Wi9���6}���q(��E4���3�(�l�P$@�M?�T���З��6)J��I�ks�i�*ȣ��͑6�
�&�㽽2IZ�Y��MK��˘�/%=��O�w짤d��=�nxn�fNg����g�h�v�վ��֕%��<@��q����Z��X���Bܿa��a}�!�Z�8
h��#cW��X����>W*�1���ό:w��0�B�4mr���`�@�j]?[J������Y�.�������&)1W�:��`51c�J&^M���A�0����.�E�)���1L)�/b������L\�
:���� �I�3#�c���:��-�����ĥ�R��5L�V�!.��5�C0�P�9�X0���R���H7ܽ��1����/���|Ҏ�����L�C�����^�����0�h��H���^y������p��8�E�/��Y���Lz��5���nV��tL��6��f-�6�+�t�|����x�l���`HC����m����֫�N1�h�GF��%�Zˬ݌#Om��-p�}�%���"%�p��Pu�߃%��ɒ}�s�� _�&�� qߜ�(�G�X�?4�!chp�Z�����^��?��2+dm�R_<�A�8�\�U��Àŀ���U <�T�˛lӎ@��:ߧVlWL�=l�s�{P�#�':^�H4R�Ր�_�T�8Z�L��eD��V��s)0ÇUzq��I|�봚��N���h�S0,����U�� �õ�T9�V�J�����*��PF%�.��|��ܝV@����M��Z�%60t�[�~d)� +�,�mPDĉm�>fto�XY��~~�!�OX�]g<)�I�b�{Yq�d+{�A�U�����	�:F��{ͮ>��I���fh������2���/!� ��e�W�b��(��/47��6�:x�J���d�m�Ci��@+-S1�ReG_t�D+S���}������X/B��)w�ن!��,�+olM���8�]%E2��dA�ٺ8a/�H�N��4�f5�N2���n�u'w�nr� ڤ��(�F
��z�����c&�>�������tk�A�z�14ns���Ek%�R8�
x�-�ˁ�\Q�vsѶ� ѵŚ!�X`L��vW�O:�[��NsJ��T��uQ��e��oT�uL�\ݬ{��c�m<pc�6]�RE|l�
�y��(�:6�Z�N,�j���6B����L��kL�#������щ���IZ��W���=������c��tr&j_�N*��vj�&� p���}�̕0�n����@�`����8%�.&n�����,��̝��CH��! �!��#z��o2!�]P�T������Q$MC�H��5?m=�}�߹�[g�sħK�9�����D�:i�]��n䓚Od�,C��K�4�&N�8�&:�&�z-��ݤ���r���W�P���TA ��Y��7Ds�v!sl�O䕷�K�L莔���o�,�����u�)H.M����I4֣���v���M��эv| ��ʿ�����S����p�����ap�i`��L�Z�i{B�x�!�k���f=�24�+Xv�ߧW���\j��d��gQ��x1� �4+���ݵ�-��FO|:���3'Q��? ��L���h&!c.��61�U�����O�U�T����}���p��Nb~�V�F��
Iui�y,	iVxV�S�x�:�^uw��}'��.B�O}�NS"���H�h������P�٪���3'���p��d�X�U`�6[���E��.QJGy*�<hE��	�m�L>��A�&�L��őy��]�֍h�gy"�TDK X��<��y�$��}�e>�"���R��$���X�o�ʱR��`^g|��n�}�Ǳ��7@�NC-q�b˞�ﶮ~�H��)�]��,��yU^KV�V%�k%妨sT%:T�MF�	`0fԃ��կR`����앃B��,�]�<�1�^{��j���U_�ڧڅ���T��:b�A�U��� ���a?N��I.r�ޏ+[["�`T\5e�~N�E^Srĥ��	n�wDUX��h��G���_D�u�&�ễL���Wrī��{�ܝ��}�=�{JH�$�Y><���??ps;�FN�����K��~�-�K�N۪�>�W;U �z�����8Q�aoZ��fƽ�2�x��bݙ�'��G1W�'rE��.�_����K�.
&�b�Km���}m~�Wja����>�8���#��d�/��B�F2�E
�tx��9��l�����i_6\|�8�� A��o��Q�M �ܞCo���ƪ�\���Jp��oFV��TR%**���O5�6���e�W���|�e���h�?����x��,�:�.�]�M.ɷS��J���u?Z&��L}Uc��n�p��@����m���f�9�C1w8ql�΁e6z!���a�d��[5�:�F����fY�2f�k��.��ɀ�Y�k:<�X��0:/_|�qj9��px����10u���>LM�S�Q)M���ZX>���������z�d&v������S�BLYMWS�8���ǆw̛���b��Eගѯ��X���"�'�̈j�:��#T��og�,��i�D�c��>�5���N��y KZ��k� Q�;@{�.t�>�ѽ��Ŗ�x�́��ӹ�3�S0���r���|��G��<�{�ď��&S���@�(�c�8;-k��[. �)��UF���]W����z����N������a�0r��j;)Fv�X;�3� �|��x�?�z�?g��eT3m�lg%ր�����$�3z���L̳�ĭ�`�G�[��6O����B�l(2=�2�تod�@Q�IE6��c� ����� ۞�[�A����o\��U�L���7�g3D�:�-{3� |��lo>�%���������iͬ�rND�:q	��搱u�+��Z_22��ɉx��	��2:cD��Q��GJ�'��4e3p��S��y1�#�zBS�֋��~ J��%�I�BUa.��b���/����Ѿ�:c�2����E���+\�kq�&MHRe*zq;�w;-ݡ/^���=/
ěL���I�vo���/F90�
=�6�OZ܀�d�ǐ���t���K�I��P����DϟD��������%�|����C�;	�y���>	j�����$�L��	��,e��n�W��X�S�0ᑏOW�"���S\fb��0o �wJ���X�F9\3���z\�S���L��4~N}lz��z�F�K�!�W�Hhv&��p\�M`��*7�+P�?l�2YG �=i �����K����t�,�Q�|y���-'&`b0�u�d��$k�p���I�>�����ʯ��H��~-������J�Ơ����V �>�5i�޳(P����L?ɢ1�Z��~g�s����{�K�L�c��P1��s�BGӀS������Ae݇=���ju��G���Z���1�k��Θ�ZW1�Q��v.o�/yx�����f��+l$�av�/��[�WZ���=w1 �s�����8��_�v���2A����ر���y,ò��3�Y�K���;��r@�smi�91�		$5v�SuN@�-��e;��PǠԜ�Z �۷��d@[�	"G��Q'��YG<�/*��k/M�$�Bv:;>� �K��"�1f���_16nN�r��v_�3��ގ�;k��o����#cĔ�x6]��s��&r����xJ����RP"�=k�-�4X�1q��2T=��=������%�RT\Ѝ������I_�]">�Y�_�޽Z��r�����������kz�I �ҟn-n4e����!E����&�	�j�����w������O��) ��Ȇ骮���2D�[�����^�a\[�23e;$�.Ed"���j!�Ĝ��m�-,	�3ػ� ��/k���-=�@䝠�7���l!�~�E����_X���^Z��b2ǁ.ӯ3��1�{����HF%���>�w���ƫ<�����X���[y[�x>��Zd�����U��^��վ�Ғ>LkB(11~G��Иt"/+t�PXŢ��4r���؁��Y�B�X�~��\��a0T�!�G���O�ٛ |�p݂�� ��3��=/����l�����
����A���}�(3���W�]v
���xD�i~'-�u�5����gݼh�W�L��19k�V&��<n�������lmCȝ�l$$ߣ*1��ՉJ}Ѳ��[{G�6�dM�H�݅J1o;���E��sn=׵�r@��W�X�\�J�#l>Y��2hs�.g�!y,Q=u�C�v(���&L���1y��@����:	�9�WK����{������5D.n{��`3�.�9o��U��8�
g�憊�J�r��q?
�K��U����kr�Z(��	�=F�4��zUdn�	+�.
��:$�y����M��pg��>��=�Es ��T/fA}��-�I՚��G�W��ujt��Z?�V�8��t�z�?dFưc��V�}1����e����5�+}���o�& f=fV((m�O�A��x�
�:	TS�0	@��uT5��c|��j���9��sR_�9ӏ_��Sn,�&�=u^��vXx�>@v�P<���TU�	#��wL?˴/��C?~T�D���8X]��٣�������n�� hWJ�d�@��b��).�%_���g�0	P�s�V�%"O�739�2�
266�u����R\+G	�ƶ�a�����z�h
O�╗+��- g��j'�9�@�߇!6ʞ�$�87K�h�Q�<)�z��b������(�|�K����"����������}#��lg��b��A\�>�u�?������u��b5�Yi�6���e����݉��6G����;��?۝��xi �V��RNR� �c8".��ݥG���y���������
!��`i�`Փ�d
��߅^��+��t���ca��CY y���	�~F�P�W��:B��XQ/�j=��Ɋ�q�ey��.�QKj����?A�'��%��;&�?G�Y�7gR"�8
��$C��3	��W��Az����]��+x��h�{���/�Ϡ0jr�jm15� 3��j�1�����;$�����WOL���4d��y��5^usK�<l�٘�P�5�a�,�M\K?����Y���XJ޹L(=��k��xV;�t���'jO�22�c,���@g
�V�F� ���ٳ�P��͇��i#1t�'
���-�GG��y�J�I�ǻ��[�M*:�d�|��'�I��� ,�',�����L	�1�lNr̨���KQW��-b�(򨎉�=#K���H}DģU�"ݗ �6��γ�\��2���'�K���h�@z�ո��~sz��.;�LG7��2�C���ACI��.e���-pU&Ǻ&�9��,c�g�M�M��#�@�tTC8��ikR�<��h��M��;��Ř}�l��*"Ϩvܼ"H�9Ý��P�I����O�i���n]#����-�o��/G��xw���XEi��1�+�h�Wlf�:ɸ����k�]�=��Gybf�0p�\Q5�I���f�
�ݚ��!uS��nE�Eml��4��g��7�,�`e�\&ʔA��j�.J�9�'	k�ϭ��_�Q~���ҥ�S��k�e��������� �e��(];+'�˵�'�F�oYe�;~�ٴ�gVM��O�4-X�Sh��x�/�,
z���T�l�<�ky�Iza�W=ILW����U�`=�IW`���]����9�8L�]E�.H�y�lm|��l�6����v�qo��&��ܷ�)qGJ[Q�g��l����5�,�5O�l˔��"Ȧd���ѣv��F�Q
c��m:��;2���P�9�����HN�b�����!��XW�5���O�p+U����<�3�F@a�!e���˼�����#�+#9�����w�N-�2�<J �_����2���:f�C;�Б�N�^=ݛD4��e�\�Z���}��"s�� `�K�7*,�G���ߡ��A�5t�J�=��5�u��D>"�;Y�'Y��!����4��1�х3@���W����싢����#�v����(�D���-DK|�]����Ö��XL@,p�+�����R�+i�Ӈ�jp�s��L������W )xA�UI���������s'BG�X�d�aY�O�;T�*`(�;N���g��* �z�1�洫L�\Z��|I���]^�g�t�;�U'�0���h��D�z�����DDDKt�l�2���Ѷ�i����<�[=B�4�|��;��quGd��V�����r�硎FeS�z�H��f}���Z	���G*r���O�(��l5C�_W�mG-��a��䅤6o��c6/���`����}<���ds��H�# �j�^#�:<�P[�t?�}0akA��D�{7�����8p�H
/��Jr~g#��`~v�G�a|�XY�?�V��c��6У ��v�Y�!�EF\��_�G�����B��>�	O�#��O����X�f��sV�0��B1��Lwު�g��z����F�x�j�q���닯��il=�?��d�.c���O��3��XyNQ�T��3Z��^2ö�H�>z�
�2$�`�E	�@5��D�u�Z����Z�ϕ)��}����j
Wk%/Z�S���F֊0K��P��ܩ�M̉�k`���C�![nM��2�R=qy�v�&���VN��:�6K��8n�^�G
��k6�5`�2<H>E��d?�Ч�Ι;�4,7?�
��@�Ԕs��=���ʅR��=�aV��������-{JOwr�e�\M:K4��ܒB��箫o�!�7S,��Ռ��5JȤ�4Ŷ*h���pN���n?w�&�m�|�p*0�pZ0�FwU5~�w��췌KJ��k���i���B=W/�HX#G$n�z4��X��88�I)�&@���i��y ���D�Ei��H��r7E��K�h�6)����95�B_E3!.�r�˜ht�bõ:�1!��q��Q��}�����i���w7��������S�C��p�pR��	U�����	�����{v�n^wO��
���l����ߥ�@������bm�)g���������xo*ޅ����{�jg!#~���D��{��MA�L>��1	�Ud��kGQ���ۇe!G����\A���z���l=��ݘ�f��?�>����9A�AR�؎����s3�R$�F����'\�=�PPHqnV����L\o���;2��m��!b�;Ӄ��Z�Щ$�t��<��%�8��rPQ�+m �ʵvOf����]�� X�dW̻P>A���>�X��
�h��������s���d @�ˇ	K�&k��!y
2��Ƨ����$C���0  u�fN����S?cb2��Ā���F^���:qqf����yx	#��n��L��"tZ�����m�-���3~b�T5ڍ��jJH��g����t�8$I[�%��Q���W��{�N�F���bf��΂�fғ2_��p��x������ONP� ����pYKe�ڐ��&�
��>�{p�6���*�g ҦA�f<�Y)���4��{<�&{i�Vd�h!p9��Q6�G{VY��] ��=�L�t%4�F�Zd.�K
}:��y����U�*�N��f��up�ИD����.WH�wi�mj�1^.�I��R���#%63�C4�B&���X< �yI(	+�,X�����#�7�ͿUi��̀��S6���� ̉/���_k��~�Bm�a���,a�`�v��L����.�����2:_�"%h�
��+c������_v/����>F�1ui26�a�u�֢����}���4S�x̵Y��)y�%���RY�'k���C3sd�rq����˭#��HmO����]Q�9�-q��ӣ����4�g]���z��g?KC�}��V"�9��׉��B+Ic��z��s�f�8�5����'����%2�����>.��^Y���|`% `�u42	u_�n8�*��.{|;O�La]�9J��}��>��_���j�Hp<��
�����O���3�!����8@�����f��t�>!����T��ԑ���E0
~��v ���~Ks�"
���#�2�*V/��eHW�L�\� ��[�0��ck�w6������sx�"�"�����G���g�v�Ms��$ˠ���gݞ{Lu�^���F�o2���p�W�Yׇ�+�Cb��ǟ�4�M��k��p���0Bo�
{��!�4�G2%QuW�'N���KŖ@O��ZT0�Qgw=��mT��Ft��\P�hݍ%�Z>J�)��x�/��jp`������a�\Ec__�m�����~:+���i�\H��/"�]u�� �*OW)�`�w��¿(��N�0�\d�f����R�Ř>"�%1Qx��/�IB嚨��2�&�3���O���R��2$6��mZ9W0����+-r��|�)�ѸP|���A̘ Ԓt��"n�Z�p:c#y:���=`z���݊�#�S#�"��C�mp� uYQLO��L����y�n���}��	�o�)�*h�/>�@��/�跠J�|$��@���y\vN��:�\�G�����eM�L�n��e��ެ�X�#xn��	�	GCj	��q/
Wa��nz6�'dP���$�	�sR��s��+��o�r��BP�t�<"�'tb<b�飬�W���X����H�������z�:0G/����/�y�
A�C@���~U�9�2�����t<��]�?3ڱ�S�B���"��b� �o��q��R�t�]�����g+w��\!��ItВ
:�gt-`��b7
��J,J\��&���(C���q��B�-I��V�M���J��X݌������@l㒅Z	�'���t�9`�3�X����=a�`30��dD�[ٛ��Ģ�;�����T
1��{3��2�(W6f�'m�2�0bk�� ���u6c���VJ�j�z�)֚��<��[�.����d���<Zx�1��YxB*�D�D�X�cY���-(Q�7�]����v�:�TV�6�y�Y�r�.�)�`-�.t�Az��V�8:�k��|����@k��;OSw����];x��LJ���#M�����I��K��N�/ObpJC��ge�Y`.| �"��*�r��qqFƊ �w���;ս�o3�3�[��6��PB8���{�u�;�|�
��t/�x<��t572iHo��?��;��n�M�F������AE5Mi��P������S�~��Uf�Կ�-��M����OP�_#oV�C��������l������O	�d�`Vt7'A���&�#|�a+#Xi�x�_'���&�ڒ$���c#�<i�����z���C�<���!	'���ߒвp��ŉ�&ߙ�9(���X���0��Vu���.�\��$a��ȼFusy�NZ���;̯5r�0z"N*�4r6\$Ơز%7���.��M>o�����+��P�)����89��j����F"b$5�۹x�eS�e�d]˙NX���Ҙ��ݰ�x�t�����8QP��+�j�����������9M��_lڐ�G���I��ۡ�L{��Ͷ�,���LB;����Z��Q���! �``P��n\��k>�iGi<��HG'/��_2H�Rh�K��3��f��oo��e���hK�P������X�e(	(5>�k-�̇���������LF
|���Z@?�x��`w��u�������_�vw
�4�rc�8�b�{���[�Ϝ�`�X)�J�w�۵@�Ć�~_��	���g��Y/1믣��b�8Q��� 7K�.�%y�Μl�_��>%(��|?៏$_,uE(z�����%Q��B����1?��8ݩ�b�DJ_fyc�tz�W+AH4�#�{ұڟ]�x"2�g�|vX�D���ɮΐ����A6˅*�$��q��(��bK�2l_�A�^xZ�������j����;�An���HTҧ������pH��2�%{ ��|�<��V��ɇ2�j��\F��P8�R�=Wԍ��P��ȳ����]�Y��c��	��[����8��ХR�J��_CV�R�L�%��A�=�����y� �Mj�=���p�c:|��r��̽�����v����3o'��ZQ�����i0	��͆�Ͷk�+����'@�t��I=�Z�)��r�+<�r�)f���e9�h��X*�Hr����G��^M���l���N��Lm����S�%���bV0#Y���|�9A>^�0�.�$-��4�"���+��!G�ѷ4|j��>� �)��n�87��Ҋ<�栃�5'���o
i��@p߇��o�~#��s�m�2��g��-ss�.~2Rӆ�\�?��{��,��5k���֍1���ӄ�bbPC��oa.K�êm�y�e\�²�f�5��Jw��k_�NZ94�S`5�Ѹ��#�*iNGת$����E;���!��O��ݢN�/�xWL@�ߏ
٩�91}Fd5�6��x��0\ެ�3��'S[�w�[W��d�Gmn��>;���������1+�+.��|������G��Kpp�=(�oPʣ�:�'�scT~m+�s�#��>JZW���k�T�!��x�,�	��M��D�K��X1���ی�j{����
#��FJ����%# �=v_�!�<nRyEN�K5S�V;��(��|]���zت�1Co�,ɰV�B޵q�\颂;n��չ^$A���(;���?����n�EN�����*�������G[:�-ZX'ĚB+k��g����н���[����sB�Kc���b����׫ʎ^�����;�t%�)"Wl8, ��T'h(5�{���	���%�N ���V����F�.7���a���XLh�����Gf;�..M�|�v��(�{DyT���ȝ_�d����~�BZօ�%��Ø^��<�~�3$�\�XֹB��Ǭ��S+.��"o�nw��.EU�I��$��έ�r_s�/-��¤�)���Y�.t_@��v
��]���y||t��SnY��{���U�	��V-a�8���j�<��u�kn��e8u 6n}T䴮��6�R.�[���e��)5���6�;s���i9�[�#�͐�����}��N3�Qo�<M�o�n�͸���y5���ӝ>4����c<��91�:��c�<�\�	~����*��jyw.�2����~t�H, ��2#��K���ikX\��#A��RĭdDa�y���Ϳ@�Sx��J�*u�Z�+8��!��H������ �����	YS!���J���IE�_�s���!���p�l��$�LI2�-�:uE�A޿6B��3��F�|�@[�-��0z�ݬ�_kL����d����)ٚ�+8�c_��H�\if>q����w�!{�~��6%$:@`|/K�e6�mNE�il Y���z,�(m�*�W^[���L�N���=u�=�a{��P�qT5�q����:�fqA��W��8�\i�X��UPa�qW0a�:dD/D���VvصT���ٯ쫴��	�us�e��;�?��/�A��C+l��w�ǣik�\d���>��K�r�:���Po�"��١��h��Gۓu���S�)l�y\T��1!�l$<�К��E�����1�<�`�]���Õ��*�2���m��Y�=:�tr��0�P�Bn��,���Q��=��j������p�d�\��;�o�-k%- ���>(���<�섦)�IqQ�/��~�1��W�����_Â��j������t�ꌥ9�ML��8���S�L��⯻��]��tQ�R��:ϼArr5!��5�\&$�q�+3�'���'kxϸnY�`���I�a�%_
4բG�;����Ee^-+-�BX4�ٜu���v������VW���ݡc_~�$���N��{�����6J�#����#�7H��c���G{~��D�Q3~$��iP��ׅ����VHaq�^�Xю�+"F�JL�.*�����yN�yX`�s��wlvMMs��z���^�ƍ�M������-�6���"-��G�4�S�Jք����(:��,��a�>��gQѬ��Pԅ�MY�1����V��թR�op�k����E��ՋPU�~xܱ��׷�g"�ϔ.>�ml墠�Y�<6�ӯ�ʦ�Y��rg0��iQ����${�VF4f\��0�H�:Qhi�έ��k?W��O�������~nT3�R[D�/;R�4�j����L�{5�s�����ŘB�|��Q���d�VW_�
��!���2������N[_R���9��9�x
�t��#A��=�j�l;��okbK�� uX9�(ʫ�s�k�7f2��ځ[Uj;Y�J˝_-��"����n�ʜ�<6����b�Cf91V�/���:�z��r���������A, 1ęGD�_QtG-��e
�5/rv��|De䥈�NAYF4J4� m����V��]dRA�Y���a}؞�.��I�X��(-Ld"��+I�GvEs��Y�K�Q^|�*��0ҹ\O�;�@�Ș��y���u���N����]��_e�[�R���Ė��=���_nE��+$fJ{� $~�ـn%Z�ՉV/�o�tW;gS�ߝ�k��Np��+	��w�j�r��$Ő���Ț�8WAﯯ�e��1L_����FdVLث&|�~�k�ʱ�x�r^w��p��<̊���X?";K�xa�I�54͍ީ
R�d�P"�����mt�i��^�v�v�����s�F�	�h���Id_�]�4.�`��d,LN�=V#�@�����cz���7�I��X<������۬M[�|��u9wu��T-����?5d�]�	Vz5x���k�[.�s�Wۿ��Y�)�z\gP�o�	��2�a�.�3���l��
��� @K�+�� ������÷��"bg���������w� =k?m����؊��ڈ"�5����xm��}�4xݕ�3�2��]�h[+&U�U,ۮ�sS�Ԑ$�:���a�}��8�W��a[��R�z��6h�E�Z�d�8[=<�p�p�g�ۃ���}�q](63B[P�ʍ�w*!Gp�	�N���� wD����]�.��ut����<����<�9�8R��88S�j�(H��,���w��@���=@��v��[�`���t�[]&Bl�����*0����׏�؀$����u��)k�b��g�~��&���΁�S�r%�hVa9�2]�6q��RL"��#�3�	S���6��'.�z��Me?ߜ�C��3@����]f�krժ;�He��vˁ�؈yzȐL��+�+�O �����ٖ��V"�C����^�>�)��޹ �n�ɁD&WO�����Q�t���@��������ل�K����G@��v5(~T��Xu�S7Gn�0�Ie�p�8"V+�]3��6u�hG�ߧ�v�$*�d)//2�X���^H\)G���oUW���v
��<��:�Sq�C���t�5zeX�E���f-����04���VLC?���gv�R��!�����wK�wݼ��p��d�?��%���&!m�����`#\kAX�?-�D�����]o���x^�Zo��(k�(s#���l�6_�&[��HZahqcl"<i�`�Y�S~�u�����N� ',Z��QeFwO�A>�5�.}�����M=`i����*�w�����$U��[��=4�mB��xvK��;�1����ٰ�_�m-���DJ'F.���f&,"O`R<)� �Mݷx�ڼ�=t`�bL�w�J�ue$S��t��e���������A�WG��^T����!���/nI��j{]�"ЈSq�4Dg -(ʬ��D��謟2Ik r���ƪ��݂����?����r�4���΅9��Fzo`�؟��`���"f���v����.�g�->0ʲ��R����sǌ[���:f.�|_6B�=�z�;Q�8�~kۛ��ځU�S0:�[�쭴�cn<�c�v��a�j����H=}�Z����BS�˅z�v$!�ռtC��(���� Ҏ��q(0t��K�c�xP�#[,牳6�R�ԴW�7Qȱvػ�u?�	�{��S���_�;1T���-���o��O��
�������V`�\��ҕD�f��ЙV���)���>�O� 	�_g�x;�R�<s�ӇF)cVz���6��v�6~UR+ ,�u0uo!P���{�M4���Ě�Yڐ�0:��� ⶶ���C���#��!J�K��E���fE�}�1���sXW�����c�34�Ry�K��˵�wץ����^I�bd^Ar����x8���*�e�����Hh� Q˴�&!� ��V'��Q�l)t�3�6����C����$��LpN��w��1_����p��(��0,Go���(� �Z�U��x,Ocy0��I��&���Ǌ��b8��"I�k���^�a��a��u�ӭ���䜸�N��k��>�i,k����>K`�DS��K�ߤ�6d B�i^H"1��>4@5+��~�Y�B����IE�%�F�}��y��DE9q-}֙�I�@�0�&������%-3�5Nq{O��MxS=�4.gu�_��Br5���ON�i�|�N���쉱KΔ��W��.#�٤�sؤP9�
��w-�Uy"K5�[W�l&�+��;"iqR���V�,]�z�1���5q(��O��Q
6M�"�$`��KD�N;�~�ܰ���Xcڲ���޾��YE$l�5f�~t������u��$5�������kAy�)�\<>5d d�\z�jFֳ�d!q�KUۉ<&�`���~��k珕ꋜy�C����{��̝��i�H�㧚��IG��JYhi��RH��i��`C*G���X>~�G"m��v�0ov�jv:���.��+@ޜ�>E�궁L���H�BM�s�Cu	m�
��oB�l;3��EX�iʻ� ������#`L��;�Ȑh���ݬzP #΄՟�<�P���W'��x��/�4k~ϣ��W��m�_-��f���z&�ONcs���j�?td�R�֜:���j�OH `��diL�Q� T"�v�D-H�Bc~!��
^��4	��۬�AOW[��m
�����9[��E7BPc��ts伴��=f�@�8���qn�ᴈ��V� u�!jI@w7�-��v�t��k��1�o�ܔY~�[
�$j<�I|���?Wm	�.0��������P��Y_�`�#a&������7��r�J���:ˉx�P��9ȓ�x�����uDć���Ky�b#݃8i �Dj�v�A�)"�s�ű�*.Re��6'$qA�{
=v�#��n$�7��}��i6�Z�_X�x�-CC���O3b/*�o���49T+��a����)k�q<��;C9-D�9�yG)�.N$?���i��ACQ��Ҥ���ϼ���uqI
KJ��k�HF�R���I|�u� ��2e��s)G�aAY�����얨�����$���1+bS���	��]VY�޸�:B������f)���Q��P��\1��c8m��9CMԷ�t՟cΦ;�Elb���&�%��QZ^�޶�Y;W�7`��H+Q���3�e�B��\�����ܚ�v0�mN6B���T/x#�2iD?\���\u�z���-�^���<���b3�T�c�s����qEpь@�0\�g��}Ǹ�