��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�\a��YV4�|�2�xrg���������,<�?�{���Ԁ�h���<&��ػ��^�@�}��ǉP8�ow3TO�-�.>�{�
q�]YA-AG����B�p�,�B�#���l,sFߕ�r1���I\� ��,R���\<X���"�����B����ɷa�c
x�����W\����>!��y�2��,#1��h�;�'a�[%���8��=#��?�^��g�=�G��a�rw��yq��+-!+#sC%�ʕ���aY���������_N�ʡ���+7G���KJi�:����_�� ���{�'���4���k˳�I�5�:h��A�T��H��C�ݎ��$
��o�Nl,�����:���Q^�Н�g�PKB�Ġ�������Q�g �*y���p�qc��p/��;o��n��h�%�AH<i%�E�kC�a�8�`F�G�$GK���� ��L���+��ث$��*m���ɀ8�F<����Y,j�Ȟ<��[����N�Q�:�������K�p����I%4�ґ������Ee�]���R����s�����K�᭿��L�*��irիJ��,x� ��V����uӂ6��ב�v�bj_
��?V9����d<މ��r)�65��X,�'�t��1C� �!�Y/l$)ͦ�ϗYK�b�\o�� ���{��ڍF�
����`�6l?=ɓ�<�v}�ͨ�n�b����#�6E2�K�F�ΜQ� �>�y ������Wġ�̴3x�֛7��Bc�jxsw��#�A2k��@�_���j%jA�����,�.�-4K˹d��@�N��������E�ťx�u�"]�0�#y����g��ȵ� R8���/�]\�<�hmג�6�S[��zo�х��,FP����6kDsߞĮ�K2F�ΡNT���2I5�	���D��k�98��$i��F���<C\V��$ɿvk��׷�9J4nso
���Y}:�������W��5\�I_j����:����~�w�	�:b������6�V��HF`U���ĩ��Q1�9��7��ݕ`��'g�q��;�W��}Z��/"G0���3ƶ�_Ƈ��A��(2Uө�
ZZ?^�wo�(Ke�C������
�.r���Az��l]� �
A��n�5�᣽FUB�KX`�߄��!�� �@��v������ɪ��Y�����)}ۺ�A�C��rB��h�i¢��t��fqZǍ�~Ϋ����|��yma)�0���ݢ�A�#�nHt��_R�	W�o�7`ޔ-A��!������n�-�xV���Hc�pP�Vqyc� G
��q��!M�@`�i=�g@�c)t����gh�Q���q�'�����	Q�/Dg��z[LhP�ی�4�&��J���Ь&�N�E����~f��V��l3��:Й�'{qٍ?,���o�>�T���_�OLB�������ܑ����{�󛶊����+��L �OD]y�Qۻ��@�zp
i�������>�&s�9�_��c;pДL�Ǘ f�]F��e�A/�Q��v�����%��^%�nzI��
����9�¿�=)�K�*s�}��"�n���X���O�B��n�U�b�w�m0= ��S������]�� !)]�2����b��ndT��6#�gr��Cmf�)�6[9�^mp��:��_EJ�Z�����3t����A[$�°\��7s���
��v�΃���Mؖ!����!�q��W'�"U�W�&���6����>=��BSLY��L+���Z��֡��|qu��{��Lj;��/2���؇�ao^@U�?0����X�W~F����[F,W�8�ȁ?�&�2�3>����x��$N����O���f���CMZ����`���.���iVX�I��i�K{0���z�%ڂ+ZO1��^}Xj�r���� �
����Bf8T�ԬM'��>k@�:�_NfM���a.W�������n��(���X��Ĩ#�L @ޠ|�ƣ�q�fr��ts't�f3 j��49�V3i7ٱ��#�p����.�|�&�φ�L~���r�f��,�N����V?n����x}!̒�.��Vf�qP>TQ��Y��Q��tS��������=2��$����tx �+� �U�6�_�G�f�+�G|����/A�f�һ��;�=&�ms�;g��^����î������f�fsVz�Gd�l�A�>�`�(l���6
P೚�!��뻸��[kS�̕��ž�+��gf� �s1Q'�)��U�1�ExJ��6��!G��
��3~[%ᅞ s)�X�&�d;�M��Nf�Z�d��;�n?F]&w�.�ˍ������.�$Z�x�U��4\]������7������qq���۸�ϫ3+U@���Sm3��
��+Q@����9�yi1lp�u�q��,4�ty�v���f��>�����J�#%~��ǁ����yĥ��9�`��'�:�^�����eYʇ兰�O�������y����BH��"K��Mq>�2��i�G�{��4��;�!v�]0�E����f����7�O���Y���|�b��p6�(׈UK,vD?�U���v�6�w��ߞ�>�I���c���,m"�W��y~%��PU��|8�Z�+�X���sk2��ۀm��s7vbB����R�!_E�����PF��m5@4�+����T�]�u��a�nP��q$<N���G������AsS�ѿ���M�:܌֎[A0B,��Tې��]9w	"�n�?H���Z;�������b����"��˂�ݷ��S�wҀ+o�j�o=���3��w���F �/�hv�0;����=��Kc�zT(��V�x��Q����ϑ��.o:�m�.�ټ9���|�`��8L,�v(@���ALmř�GK=�'Ѷ�n���,��re[�9���Z�N��e��H<����Z1J��[ڳ=�я�'�09]��Rqi��9g��'/fj� y���6�N�H��u�1�2�n�Hj�b�-g{��d-��Y�<�t��jx;4+z$���PJ���L���)��dT9��ѣ�s���^��"Ň���{U�QYr��-ڳo�y)<�o���A���ʩ�����%�a.�켶|�2QD�)@E�K�����-���3*o0�~�D5��S���E�ܙE8���6٭���.K~���jբ���1�E4("��I����������-z�����*j����	;9��A���%G�Y�N��I��ry�"��|4�\X����Zd�FE����%��6l$��ě�]��}<i.,��'��|@f4����%��Y��������=��X����=y_��z��_��=��=��eO9,f�9�h�k U�p�)#1V��<�y�����j��y�Y�ˋq����h����4":���f<g��Q`&m@� ��KB8�~9�B������;�]͠�$b.����z�����@/���q
TG]��8�(�1?�eo���]{���
��:\�����6�_�?��u4i(��_�� %��m(SL���Q��ϗ�T/<��\�{���`��Ӏ��>7d�|^�N�W*
$���<���ȳԤ���Ѣ'�po%M�)U7�vG�>��~���ԡen��cے {7�7���`���h�y(M4d	��e�1��e'�s�fo��#��~N��� q
o�v��� O�ȡv� �чR�Ƞ��3��G�N����фa����B�u��*�Ez����c������S��������e���2h@��J3	���8f���K�r�RZ�>�M��O$��qJuhn[���Z�b}��'�֟��0�rg��2"c�S���V��_�x^qp��4vo�nA�<jh�&#�N=��ˣh�d�s��Т)�)��uS�ϔ@�����l�ͬ��Q��i�SR��"@a������ �ߵ5v���(����k�K�KE2�i�e"RRN�x¯w޺������V���]Tj�z�C��I���̵-���-񕙐��8�����O��H����|��l�X5T�`aG���lRC���.���	�+�3HQ.ˍ#�F��e�6�#o���Ո6��^6���3��:����j�t�颵���0�:�ne���݂��k��&�o�����{����J����{��1sbN1�Z��-�8�ua�J�	�+��m�/����9�zw����##�O�9� ��@��"�����=�g�)28tȊ�+j���C��԰f!�c�;
0qa��� �����-�c�N�ey&��+*�&�Se"P���
MWt��24���p���$��Y�� �{^��ۙif���W3=�/��T��,+�� ٰ@���D%�z�����U��s��������������q�<�M�w�G���6z���:��M��J`���-%l�?k��x�:U�dBq�`~X��`�@ �Bۃ竍�q	�"��f��N��F�.�a��=��w�b�7-��6�)"+�+R�5�/Xχ���3_�l��ڌ&>C9�h��@ˉ4RfxO����غ'>�_3��LK����Eu�ą�͞�*���(��`��^&uQݞ/x���go����ڈ!��CE���pe4ܨ���6��nF@�@A^t�o�\�1,z����a�(:?�㲊��qG/k�\�����ngM^��T�s�W���oW��a�nZbԈ���Y�!q�L?��CZO�<��|��ڏ��J��$]q;ߐzD/�-�&��a)X���i����2��f�4���=����hj���,Jԅ�m�rFgtձ�B�W�Q͕� v�[B��'ۻ?��H�
�"�g�8�6�L���a��M�)��B������r�����̮��9�I���Ǧ����#F��	@�18�xbJ6�e���0�C���c��>H�l/��~1H���/�\�3����p�}���U���C'�&H�	�y�.ǯMk�T�0�e�'E�*��3��I .9�����wb|���q����ޢSnW�tǢ�q��b�
e��Id�<�G��!:I�cC4����i�\�$��[����$
�O�<>��$�5c^�ۚ�i�l���}��TH�)��y~���	GZZ��r}v��l*����e[�Ig���ۚ)���Dd����*��[����9�����F
�]��ټ��훛6��4��IP^ۆ�=������u�/Qj+��ѳY3�lo�E��iw�^s�h{w��t���t.ʶ&K"�m8F�v|q��uau�2��J�`��/.t���#:w�N����t�4_KI�A�֞����W�C��2;����E���K'�0��wg��Q�|R`]�!נp���RAȪ
��:�A����Ә���w�.��U�L»ݎ��{$��F��Ixvo��p�lKU�8Xj�����vl&Q�$f"�ϧ����WU%\=x����P�OH���qoN��j���x�����=����K�G+&�Uù��s���_�_T�E�M��,	Jl =��"T!�%oMz�?�]Bl��\Zfh�j��)������% �b���vEM�?6��:U�+�~zc�����ॆx6z��v�~��?�������.?�}j�ca�.`��W�h8D �Յr�|����K��j!SyX}�^P���L�	6�z�&:b�n�q����v�B��(7uƛŇ��Cp~��/)@66�j�BV�� �r+��		Gb$�Sz�x6�:d�?�������:-W���i�:��Y�C�2����k1!�@�N$Q��=~���ߠ
P���	]��MIHX{_���e�\�Sgw-"s��C��@GxO�,�X���\ޞ^��f� �������ڎ�ѓalgί�7��5��G��	#����M���[��1#��(����	�+tډZB�>I�UH�Fjhy7�S����Dq�i)}쏦o�`Y+������LS"�� �\��'��@z�NF!�tu��u(�0�E|瘮Z3��tL����ü�<(F�u�����a��P�!"[RB$���X�C ���5�:24;�#����*OF����G��I�}��#����Y�vh�35����c7n�����\Yd�J�rQ���>��a[�1�z�v��)���_0���x��ӹ��_�bkݸsƬG�fSn-?��ۢ�Q�	�7�W� W�敽�v_4fQ}�ٶ�٤yb��^cq�	_��RP<C"k�-��J�%��>���(�T洭��ҶO1C[s5�b#�Л|���XK@�6;��t��v��Ơ�@��=OP'K����C���0�Z�w=N��Z��-)����f�j�'�j����.@������:�����´�z3���Nv��wndR:�Fmc��}�l�Z��\B!�G�6�'iɚ�9�e�D��}uR��%�7�b�\2��s�(<j_X�jf�z�>��s�bqꔞ�aW�.7)����
�iEZQ�����@��J{��Z�4�^���u�c�ˬ���4)��b<L����R}Z��9�rn��3�`<�8E!@����1���ѝ�N�"j�ų�>B���-�5A�����4+���%7��$��&��J})�Ǘ���V�k�c�SO�ub�aDT�p6lZ���{�F��5���<��Tv�~ɂW~ǖ��V��U���B��sRv�y ��Vxp%��}����P�싪��+�DV;���"p�4	U��0�?K/�(�s(�e����=���U�����o�du��-W�^����=Y�n4�Lu���{���S4��Zv��g.�A�;
�ϣ���|�to����+�Zcul��VP������2Ļz%�1��k�f�|��� �������Y�8V�P�[��g�q���>YaX/�uC�y��Pf����lqA�8 I��-<���]��� ��c(�����	�Y�E%�� +���#C�uk_fb�������Q���F�-C�(7�V�p<�`/^����DU�\|�o��]�F쒨����P�rS��F�p��o_�5TW�#���x�?�%�j;6k[�ScA	����A�5��ʎ�����9G�B̑�=��k$����y������l���8�JO|ۊ��!��g� w�Z��B��5�ݚ	[nП��e���8܉ы���˺�J��f'*.:��5�סVa�h?��#0�K��9�#t8�����P_;_�m���m��Wb����:rb�ȓ�z�Rˊ��X�����rH����Z�ŕS�B������Z�ԫd>`���G������>29�>��Vx�)��n8�И1�6Wh��G+��G��$��693u�(,�O1���^�^���#�w�ux��׺A�ȁ:�8�؀Vx�"��y��v�tW67q�!H>���lzD��<�#���<-�W�f�3~]���0�g�f�d��n#�\��ejDtOq���;�E#*&�	o~�*]�{͒�/�_e��s�uF�5t: ���
{:��H:�����j���A=pP��k�)-�9��|H\�L����z$)�I��?�������cՌN�)�����̙7��Ck=7`+�a�׍fE4�����5l�5sa���4%��aEg�o�2G#>���Z:˅��Y��h���yC��'�fs�j-�����:l�υ��+>�㉻zMGyl`�����9�|r�¸!-�����_v�p���#;c�v�,���<0�Zo��\����'1uw;��.��d ��σ�c`[s���QMC8�����K�!ܕC֏��,�OЊ,�fYMn�p^m��]���Gg�8���gB�L��,%	�LȽ3v&�!#�O����c�K��|�ǜ�Q[{q��7�5�Y	6�Ê��������Y�V������Q	���V6� 2U`��V���T;ض�ȸu>R�8k�k��9�7��� @]�L3ܬ�R���Z}a�[n����3Ö��
0���v8����hn��6�����>1��h�{�.e^��`��őH�q�\.���EX���s|��k�vr��̶�䒦&O`-=q�P��*�p(���j�O#�*��'�GH��D��E��x�l���lS=���Ǻ�1�,�:9Z
�8R�ݢ���G~A{7{5���.ټ}LƟ��i��B��_	6��"±�dZr&����]������@M^[��K�C�����A�M+<T^�`��J=&l赆�S��ٻ��n���w����s$�	w��v����H^��!��י_�����>4��'�>�/�'��!�&���tܣ������Z�/bbG[���st�q̾>��~��evr����&�r��	��/��?����]���Oi�\O��4���T�|`h�	�� u��X��;j�P2�{��\�U7S��F����;O�$�d�A��i[�lpB8ٟ���k�vGߌۀ9�O �G�ϰ��(�M�~7�����}۵�� &��< �l��ϼ����]�\�|)�vm$	�غ��'���%�`�&�;{��?#��y���!�A��x�p�$��VB����`��/�æ��v�_��"��O{�7�uKv��s���f�N���?b�+���ĵ2�#����^�����A�����o(GAM��%͜�HĐ�VÑ#�ȍu�0�~��q�N}j���);��jf�#D���k=�34�|��bV�evt��~���+�\�@V�fHk<d��"�FɄ��SM�A�Z��l~��>�
O�W$����ؙ���4p0]�<kC�ݬH��BtȮH�6hǥ��VK�Hjڢӯr`_�Y4���A��mn����c�d_�Yڴ\��$�m��L����y:>JA�\ߓ�@c��%�j�px�O��T����t>]�2	hT�W�Q�@���,Z? �n����i�C��q�����h�^��](K�:�6��Qɴ���B�
b��[;��3�U��5}E�����"������c=�}��Q����8�ߙ)���L��T��c�! ,C�Vi��Yœwm>4�Vr]oB�� �ߢ�9�
dϐ^��������ֶ�'ӝ��3t#J����R�85�h4�	��*u.��z����r���Un�"�7*�}G�d���;Ĕ`P�!�Î�Bsn$0R����J]�Yٟ?�$OL�ǳM��WL�Ɉِ���d	�W�S����Z���׍�2.�v��PgZ��&��+f3*��|Oh�ǵQT\��J���s&�=/��ۆp-�l!��x=��N�ݫ^%z'x�ri_>��>" ��f̩�|]��PscG��&��Tz?x������/���B�i�Xn��.v&"B�0��[���p�b��(�b$QK?�*K�6w�x�ﯢ�O��Ҵ.I��^��s�7����X׻����<E�G(���`��֖�D N�ʚ�\|�*L8H�r��#��������<b��^��YF�dx| N��ܩ@n�g�~���� �F�\gWY�6`Y��G$^r����AZ�c0��%�_ү҉����	xv7�ȡūV햟 �g��{���f��^=O�xl��nԾ�^>JW-�5|\�ފ��~,��*ӽ�u�k8D����֛ *3L���p�����'�I�F����v���}�wF��h�J��x})=���SԶ��>ĝ�gCt5���(3��.{�S^���_�5���)Pډ�q*�����:[�H�q�P��RY�iB9�H�m^cS�E.����\9):����=��T�r�%N����	����#�|�qq�.ѯ$�bk���?���ǅ7�,p�����%�4蜤������	�("�@�aZ�-@*10B��ȼ�h>)t]� %�\N�A>�$Zw�7	Yh3��L���Y�� ��a�G?\����}}�eZ��PiW4�6�=��lE����e~w�Fʝ���uJMZ��`Z�ʯ,s�<]ܧ��H9��YW�|[҅j�xԸk�?�7��u g	��1��g�젼�
([��_��D�)�<�n��)i%A<G~>WmMٵt�����"�`�lʷsD��1��y�a_�G�TE�N�Y�k�{�L/*�,e?���<��B49�?���/��L+t�^����