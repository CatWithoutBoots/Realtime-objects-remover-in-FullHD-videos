��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&��^L�h�m��uXҰ)B��I=��N���f����5
O�a��Yl�Eج}�DM�����,�����ԋBQa���R
f܏��)��d��;	0d�:�1���t%)w��0�<aR��ք��,٬m-ǹ+������x�B:���X��9bє����X\E'X$7�w?&ٷD��w������&�RE=��u�bJ��G:����������UƎ*�Ѷ�|����&�ie��#�6�u��/gw�L皵�،Q;�MX���Hײ�G��pca�)i��z�'�'}�x��J�p�0|�eP�"�";�K����cm#��UTG�x���.�?�D�_IC��^Ɂr�/l���ǟwc��J������i0d:���[��/Z�9f��'���Qȼ�¡�E�¨_�����ŵ��Γ8*܇=�<���P�[mOӠ�5� �S&��[��k��8����ž�i?F��c�" )5�Q�����
���>�xF��NΔ�e�r�,�i���g�`i��k?��H�Yw�+����	G�h�(j7w{	|��?d��&(���IN _<��^Z��� ���8Q!͓h���'9���(l��E��[�|��
um���Zc�,��嘑��+lC��yÞT�L�,0��⮲�T.�m��wKYtѯJ2���95.�sNyM�4�Fʲ3E��2���=iBY{����.y����������[~p,���SWi^��WN���W�nn�Q�(�q�y��;T5bf���DB��8�AEv�/\J�6�fi_�'Y��SU)z���>�.�f]i��	��=nX_���Qʯ��^]aN5�d%�Fk�g�j��R���hZ}4��3Ӟ�+(����kkt�Ƴ�8%�̻�ۙ+�p�[2��W����U=�1.��憑��~�n�i?+���R��Hן��0� �0Y��{��V��fF��he3HS7�o�����b��p�cѯ:}�1��O�Ku�{���(�Sj��)ı�W�Ǽݷ��bԮ��`Z�D�/SW�D(���ͱ����R4��r���)��F�pT(b�y�_�q��9Eq�<m�'��>�6�>\8$ǒ!� ��׾����3�MXH�ӥF�����z���7��F|��e�k$���7sȥ�z�Csp�����B ��i'Re��m�ǿ�U�ٸ�Gr��!e# �1u��J��6����XS��5ݖh�&���Hn0��
�P��8K��'&�^1SU�ۧ���2�s�Қs�̦wR���;ݧ���%Mgߎ��Ü��88�"��H�W��w�K���)F,ri
Ўρ�Bn+��lo��w�1;pa���,_��M�}����_W{j�����k�/>��;~��qa�tx��U�g
Q�h�~�xf�b�m;������(� 4zR�R�w��;�;ٵZ���>��A]�7���*B�}��?�]���~:�ŷ����ڶ�f��-�x�N6qKy2�'m���|��ɧ8���PCm]��z���Vn��VMJ�A�}��� ��53�E��,����[�آ���4��t1i�)�SzO(+zێ&�ײ(,�i�d�:��js��V%��Y�u��ir�;����6If�/u@�bh˙��9�܏��x?�~F��ϑ4ži��\�I��̏\vt�֐�Q��Cz�@W����}�M~'s�)Ζɩ�!�q����������a�b��$R�,o��kآ������SbLm'�K!��a�>Ƈ�^���'`~ϛ�vIM	In�Jב�#-R�C��7UO|+�`�h�AF�V�,��ۙ΁u�yj�=2T'c�b���� Ώ��>q0�ꭾT�����f��	̆ެxW(��J��D��Zun��B܎�9ց�>�i��[��2���/�C��H׽�Wٝ���ݞ��(=Z���~
Sb��~���í�K����4��"y��sܙ�-#�4M|�ŏ�c���i�&ϜM�r ��q~�#g�H�v�/�RC�IW*�	����� �L����L��j�����D���!-r��z���c�罎��aeLoW&�U�IO1t�_N'`p4��2#U�9Ј����򂗈S�3T�|N*���q�r��3�񿠾��<�^�]8��6g`@���]�(�cW�	V?�����2�a�Z���z��f��p�N��	E[ә���jEe���ȍ�II;\�Y6 7K�Y&�����飔
hS8s������W�פ�^/%&�uX4���8/G3����'N_��� �(]�J_.�K�qZ��.v���X* ��B�����	3�{�֮��#�׫HfxU©N9E讦n�0�o!8���"#y��ҔI��m�aӳ�ܱW˥��P��,'�k�p�Բ�1�3�u,�^�NbfYW�����BtƇ�q�eCnO�  �dN@���0��I)���N�0 �M��y�!���8��K�g1����~/�Y��p��D!.�7�[-�!;x�'�%�ś1� 6;�^�G�^�9SRx-�>�A?b�z���[���������by ����1(����;���J]���:K�_WD�k��i=�
a$��TYk�=��/6퉊!�.q�	�l�����3�d��:�-��F;�5_��&�r[���8_������缏�N��j|�w,��lc��N �El��m��z?���灒!�a ˟�Ҋ�9���(fu�~�L`8�X�L���e-q��>4�͡����s�-]��
▾K}��;ǂ��͓ro���X�ۆ�m�I�َ�"�N�F�J�P��G��6��iQ\�[M�#��ح�W����N�h&;i��)ŝyMKVя)��3�@�-i�E���$�<Xe-���hk.��)�	����%E���7�U�5����������*��g3MP���jE�V+'��6��{hl��lC)(k� xT��fI�CZ+���}ͩ�]�\&�ҫ��-a	ߨ��X��QX��	�-n�ӫM�~��c���]�^5�d��#mq�6*?���e�4�:�O5��?�n��Ȅ@.���+����ܩ��u���Y3l�	��e�<�MT��Ho��U_��Jw���2!{_�e��@�
~3;�m�0�X 4,� ������!i@�@J3rO)Ѹ����1x�Y�����%��E�n>�3��Rn�sK�ᗉ���P��tf��
��J`	x������.H1��!�Pw����u̪��I�0����};d_��=�G��K��s+����!޸5��;�����]�.���trV���j*|�-��}���A]	2]�m��y���c�q典���ش���\ ׹QN�V�s>R=|�CP�/�0_�vr a4�������R=E�,����˂V��Ĉ�}����H�y�ڊ��IU|�>0��Mq� ����J��I��nz�aq��W���	�/sn���[R�a���dWd�y�J�q�H[�ZoF?ge2��!��q��Rݡ�4��x��ϪK�1Ŏ�խ���keA+�x�o�b6�G��v��H�e<�5v�Q\�M���X%WuC;���-��2?Ƅ���ݵm��k8avX�Ob��1ΊK�|{-)5,Ъ�~�~c�:ĸ��1�F6��M�ł���Cʅ�3����������#��y]���Y-��e >�c���T������Au�@x��@~#c�Hk���6�V�I]���G@�Z������B���'][8�v��2BÇ��W�0[]4$Z��b�����1+�qKI*n�R�\���S��f�5OPU���<�S(#T��\*�O�GZ���O�[�O9nFSP�&VH�>YB���m��&��>�V�5j/����vT*�M��М�Rr"��A,���+���֬�G�>��+]Qo(��n��=+��H�R�L)�� �����|~BP���I;Re����0�q\]j�a����&�P�6dz���L��?��/Gk^ ��w�gZ���`�����X	:�ݨ��@�ez�&�a��k]W;�)a�-+��%޲�8�E��7�8,�;�`;�bM���G۬��*�^MOF�@IKkdul��4�#i�`J ��ً=ϐ[���O��@O����a������+��֤��� ?ZXȭ���:�b���yL�h�,.�D�V�T��H�
��L�6h)��x�>~K�t~@���u@{A;|��=�!��L-:̩��_p�XA��8�k<٦~�H\�v���c�{���B�<.�Or�>w5Y+���jgn��v=h1�%�l|	�)�m�,0���[v0_�O$W	!YyO�v�l�摠+���E�ֳ�_�o��W���u������C��@2���>+���7}*$#���gU�2�ͥ�W�=B���Ԏڷ��͇���m���0g��\��ř����n�K�9	���쒌��k�HT��2��R8%Sߜǂ��M�+s�5���ex�.��P�N^#P�x?l3
�:�i�����L]D!�e,)i��tǄX����,n��[�\Nz��N���L}�mF|ޠ�h��t�do��t�I�
Mh��3��B��h.*`��/��ӟ�EY������~�\�)HD�R3ygU~e~�/U��.��D<tx7��N��r��U=�����o��eX*��&/�{������߽ �>\nw34Yq�A3����f���w�7���0k:1Ѱ�.�NF�b"h*s����R'J���.�4��ےW�$�ޜ������Q���Àq����HSpCq/>lc8�#�	�V�`�d#U�"����L\4,i��N;�qS�j��_!5����n��UXH��"��-����G�������(�Oy��r�����043��6��Q2��!���meӅ�xd��j��i 1T�uâ�Q|��b+�?@ˌ�C�#�,W���fӤ�9 'G������@��=gTz�}~3���:���@�����j��&������lz��I�����(Z���9���i��_R��*�'�Z�6N���w!!K�G���+�	�G(�EF+���kh�U�	�0?����A�� �d��S��u�q\f�@�S�E���'Xׇ>���b�v/�t��[$���ms�e[�3��%��G^z��1l�&���4@��Q��7�Έ�3v��-������|�+gJS5��n�j�J]���hR=�)m/��kN�sa�[cq�.9��"�^W�F(K=#����Os&���lX�۰�-��?ԯ�\�.1�mMb��s'ͽJ*F
]i�B�X�`���C��r��p)$�	�<WO�6`�$�:�yM�H�����M�@�����E���(�L�)�s\�tդ-Ks�Sy9]�S�K��5G���S(K����r�����F�BSe�o����̏%py#��5�#MT��6���I����Dk�4��:�f$�ϐ9��'�^�8+�����C~>)k��X�xS�uf~G���0��	�e�����ÇH�W_wN�o��%�GD�!��6����`XP$w	��#c�Iu���	�4�E��P~q�t��Z��A��7�,/�f��!����%nđ%�����0E���k44���g0�^�e���� h�2���s��*�F@���t��J�`�q�T5��|�ǹ#�����?��7���9�=���mW�k��
��
�����OlIy�Z_��	��y��ET���A��=Ű�o$������G�?F�itqS����ۓ���2ƥX>]���a(z1v4�����Xaf$Y���i_Q�u�l�,��=w�qz�&�_nYp|�ں���z�1�$$��y��U9.�N!��z6R
w��^��͓�J���Yt���%O�����4HF"��z<[Ǘ��k ��S���b�gƴJa|��-���UZ]����.���+#�\�[���Tz�+(bQB(��y�~=ʢ�s��l��4�5$Z7���\�����Vo6�%3�p����=�"��FT���~�#0y��$CF��`��a^���@.��ep:!c�6��]2H��;P��׭�չ2��^y)���Y���j�������V�iU�q?���&��ŋ2D����c�'�u�����i��&	ܷ��v8�ܡKiw��pa[�V�>�;%�nsŠ)�0%����:�U�����m��[�@��t����f��Ht�Ѝ2�~��������_�	���q���Ṉ �/��{��kHr�y�ʞ��ٮ��f�eLoÿ��_V�|�un̋)2o�o���q�r��f�,&ou��t?�e�����W?]��q��/dp`E��Ig}�35;٘7x�2q���d��̈�S�L�po��R��sխ��,N٨��Rc���&�v��X'9 �u�ñ6[&ZUQ�w��g��Ik~��� �ӊo"oz�̕~�ĕ�V��6�:Q�eό�?J7@�͆n�r����<WvzM�;$)��2
�?3�y/��ͫ>ve��̹�ҝ���F`N�綧4F.��K�p�-c0�L�s��5����R�C?�gٮ�����l����P���sС��1<1�- LIX�Ϸw���4 �S���ikFkg��K�_������BH�!P�Q~�`}8���_�Tj�es�k6AϮ3���W,���ڹ��}󖬯/������@�v|�z.g�1���g�hy/�����yhcI�at3g1�,gq�O�����v���{�L~)ap{T�W�qe�0j�e�2 �n�rq�!�\grh�;�&��T�%t��c�z����{"��U�Ǖ�2w���	h�8�ٙ��x��F�,�W�{�4�|I�?�A�Y��-b�㚴ռ4��:���n1ǀ���g���Z"��'&ǅ|�_a����߶���/٦TH�.U����1����A4�7�+���
�DH�c�ɈP\õ.����vc��)�cK>�u;��+����Y����{�xdVLl�{ӂ���=�I�3�.�����]���8��#�EY0�㔹�8�@�{�#�tH���^&����I�$��SJ���3Kd��\��ʡ����S	�Bu��j���r���[�È�1�gvtя#UY%"�P2��F<V�f�[+jtв�{9i��N?'�л'�)��4�� B&�c��?&a>�(�A�E�$�\��0a]ɿ�X>�4j���/�~B�Y����7^"��I5F���>�=�3�Mt�PAbݒ�ha�YY=�Yʹ��I�'{�����	��c"�b;9Ҝ�kW�,���7��L�Y9���p��;0h��"BZCt��rc�+�3�C�9��ؐ$��*���!x�$!�Y�z���C<�쾨�x�ȡˮ���ݓ�n�������5<��$����q�h�H	����|G	cT5&젅��p+M��{�|�y?@~����h4����H���^>OM�d�H|!�Z�����ңg�A���^Y���e.�cK�o��*�D��*��nN;֘:�J��ޜ�$�#ϠA���;b���&%YE���d�u?=n�td�<�L� �H\8�]�o��M��a�;��7]y�e��L�
���rf4�%*.e	�F^�s�$kW�CX7T$�\����ԑ��{��l�uօ����T��{��e�yA�B�o��ۻ� ��b ����Q*����6��;��=ہ�9����ո��3��`����e&A&O9��@^�&Zq��I�k��z6�I�{������r(�0�4v�^�\B��h�����Pa57>j���/x�`b�z^�xEհ&�糮���F�7?ң�l�c��p̨|d-�Ė�m�A?�g�|���� � ő�=���,R��|�ԗ��uѤ'K|j\ƫ����hC\�g�Ϭ
g{(��j���Y���z�:�G����!�c�[�0BD�B/�v��م�ml�c��3���B�f)>6N���E���Z\�%�G�F0q�����[�A����[	��d �4`�cu��#�nX����o�s�c�{������U�W��)E���#Ͽ�4��I�@Y�ǐ0��{�}E�~e����O0A��Ex�B 4"�~0�7����9�</6X0�dy `'�'��F�$��miO]����?K}
w�t�����rR��0��g��'{d���Rg��<
�P�]G8~��~/"I���:��7�صM���n��"f���/]E"��2X�l���Zg̋�Dd
^�M���������GO'�X���k0�a{�\��6��t�kX5����i�U��9������OG���b;��
I��ت��h;&�bb!-�������WF������"�&1.瞥���2=i|�>^*�7�\��
�+E�� ���o��x��A�*���B>�:*[l�Zh{��jN1�N|�<P,A��š��C8@�2^�}L�(1s��g�$`ҟ�UaIi�Ӓ��j&ffC��֬�yӴ>t6���ԏ=FȢ�(���{9\lO��S� �($����N� r�Hf�p��0;����1}���(4�!�E��	�nE�q4�A����|K:��͘z;]{Tu��T�GaÆwv�qO;-�O����?u?�4���u�ڷ���8p��WU��ǞU$ҏy�R�*N;�c�-A����6�+n[Pf�,�o���1�b;�����d���T���|��\�m�:Mh��H��[˅��J8 ������䍑&����7���P+�����z=��`��6sl� 9Z�:
|�m_�Tf�y>��6S����N?�X��F��4�:ZzT�G�x5ڟ.+�!f�]'x��* ��ϩ}���kz(��ځ�0p���2�׍a�F��i��<H��R'�x'�-.��;�͹���Uq���'l��"��:�1!���5�77�b�{?��9�N�Q� 
�l8B�|������K��җ�[1S� ]�G��}M�b��f5���@���`/m[GQB�"����n�J@Kδ��]��Ւ�1=��'��.�x���|4q��Qɡ>��C
������-ȻB~Dgwf�H�u�ݟ����@�e��ү`�6w{14T>@�O�����u�Z%�M�JON�s�db�Apzb��1V���z]b e$�:������9a��?�@?�{'�t{�/��.�t�!@�ۅ���/��8AKr#t����ղ�������o؇3�<���T�֯te;%z��z����QF�w�Q��v.��;��h��r����?J)�9~O���>����b���X P�1�V1lO7�ԡީ���_�()��P���Sw[}���z @�X�5ë��"U�&8JĂ@��"j#�8�e�'��R�x0f�����
<�#{x�ly$��¤���y�㒲A�[��۾��>6zu����>���U����Nh��={ۿ�����R>Ze�\�����R�D)�����oe��!ǯ�,۾�ٸ������	�y%��n\�<��tAJ�N~c�>���^�[<���aY�>,����]@S3��O���f���mV�ģ�&�j�9-��QӶ�,���K�[%"�ޝ�ߗ�?U�p^JG�|h1J�±�R"�3��a>M�<���("��l&.	nP_Ώ�mʝL�ە���/Q��	WY{�1��fs��������I�%囈��c��%XxBUhq)u��m�yO�Km.�na�4Ɯ�n$�*T��Yt.�P�M�d��g�7[^�	���'�$���8g螤��|ؙ��HW�H!�lz��O�cF�+�C�I�X78�fs��ƿXc�|�Of,�ÖW;��pMXT�֗_(t��o�mGT2D��e�J����U"�s�bU�S�$�ƽ���;��}�:� V�"Ku�sŏg�\��d�o�W+ A{p���kɨ��m5�9��bj���0������@�nx[2�{ �Ǔ�JS=E��*��\s��T�4�f)|p8&�R�2]x�E��|�D�d�|#��;�0J����Jj�$8�>_��y��s`ty��g�:�T�BY�{D�괥���,/u��%&R���T��C�~u�d��2�y9�5Z�n��nT�i��Fd�(/��aDd^���G���ه�.?�$Y�@T���H��j��v��6YM�1��^���=��v�p�ھ�Oɹ�2i�x��\��aq��K.I�`S�<��ӕ��ne;�C'�1`<�l��)��^�J������HR�����U����y 3ӳ ��.q�wϴ���6W�9h=��k���)����F
�,Z���u�q(!��>�	�!�u �^�	ڲC�_��䌩I�{�
��dDt]1��r����]7u��I��J2�v�V�M��A�;�;�~�h-�x���#G��t��;����J����X��!f�O�~��b3% 3M�2��z�Y�k���26�Sw*20�\Ν�g�CJ��.�����#���~~���n�<(�ێdLP��R�{\�s	��y�`��
6`3�А�%�G/>f�{������8�8L�>q7aG��d���R �%�46i�
+��.�.��PV.�$���&��iq����7��w�.�R��Y�~a���K
.�yN��sU�FP��z��:��H�,��<���H�]���<@:0��$��b�G����J�`>�ʯ��˭�t�E8gBw�츒&w�^ʽ	I�w'�/b�J-F��r-�����ۢ�P�j�҈<�cX�)Q��p�e9|Wn.��[�W��1����]*m�	Y����y�6WEn�w�/���*��e��mɳ@'�B�۞������/5��.�0���4V4=��R6!=�����B�j�g֚�׏��~L�K�Mn��g�UYi%��k�ǫ@&:�t�dS�=m�����d�|�5Z o����?�ݤ�,�$
������S����1I/Ǟf�YjY��HHO��Mƶ
'Uyd���bc�H2Dw1�ħ�:ɃkW�m���X��� �rڨN#�acL��u��ߎl�������Z�����^T����>Z�>�b�0$=��D�\�s���%�aE>9G����р����ۧ[Xwl�n9@���T%m��YP�M�ȱ�2뼺��`��u�Q⟋�!d\+*���������/ޞ��N�`���P�����v((��4��ɱP�?�!��R���7���Ju�Б� I}o��H]�j?�1R���w{)��$�G��$�Ć_�ja��Y�\�ߊ�:t+�^���U��rX�R�g�j�/���Bv;Z]�n��\�G���$(v�d�ldAJ�"�$`���e� ȃo��h|9c��a9�XJҗI��ȋس��#u��o���>.vn���~9�t�)#X�C	�������o����:�J�:xݛ�
�?L<IT����<s'h��w�8���������9���ɹ|�i�5��vf���*p��;`�U�ͤ�S�0�Js(���;�1Jf/I��+lR(�� ���Qك8`:����'E��n\R�2NW��`ª&��2��1�μ+X/s��j��8s���D�:RI"F�{���'��T�$1?F&�|0�����ҵy����׈u�Bڝ,������b3���?���M�S�����!�À�5��jpH�6���$����
3�t4�8ת�E�y�߹��D��Z=����t��r0��+��3`����kL;���A�n�BH����m�	�n;�{ȶ�	!�������r�U���e �sP)kL����_�}'��vK�|�Z0����cWh%���>RY�֖
z�0�yك��S����z��Q-��N67,.��*�̣������(fO��vWC��۱]͌�<{|�D��ޡ{�(U@�&5�b��+���/b�Dj/�ָ�1���R&~Qh�h��8�8�?�.��`���b����9>3�s�L�
�?v S����]��~2��H�|my� �(��4�0G�_fXj��	(#��.��W��WZh��s9lw0y�xY_����i'�m)��t����+��LA�0�4+�i.O���\��
�}���TY�6��n��V�9pPLz�0����Q�cf���éP`�QceI��PWm����N6�%ֻ�ߕ��M��{���j�:�J���D����|N1�$��a��QJ%,��Ζ�9t�#�J(�.���ۋڱ�����,~&�֡h��\p�wrf^�=�{��Rm�-�q�y�%��ǥ���˩����L��>�;Qx����Q&�3�\�W2�ե����˩� wr�	�t�8�b��� �&#����W�%�iV�z����&��FED�pL=2�7|�:�_���U&�]P�&��a�j��n�F0l���3ƺ����vB�h�A_ժ�<�h^�;��Ӱ������zF�z,��F��HV�UuG��M�4)�FM$����8�H���|w�ƌ|&ǃ�;�I�>ba?o�1̃��Z�}���]�i���d6)2�5�Á�Ƕ\����ꉠ�pR�>�����
$>���W���,8�1�Q�{�v�³�H��k�H�Q��Zǖ�)k�Hx=Ne5}�~�ap�a�"J�(`b�� �jDY����B��p�<Fgc�O����BdV�O�{O��d*���{����|�s�3�7%��� H�Qcſe��U�S��V	:�Q��+nt) �%%�V'6�0V�p%q�F{�X��<����0�i�뒊���g��tOA�H��v�����㖷��D���%P9"9�>��=����!cُbJ|��Q$�_�m)J�� ��"j#�Bx�Zz=K��Rƒ�!q?�=Ķ�|���EN�a&۾�J�/�DI1tG�!�'��̟1�;�hs�Ƃ5��λ�Ѭm�\���i-jn�쵪˷G��;���d�� -�~"�����A�B^�ŝ�y�5��3��pùC�O�1�-��'>;�=,ŗ�1�ke�?�6a��l%T���J���8��z���ί���܎!��ز�@�Ѽp�UZ�`��ϥ���<��/E)\�Ba������A�l�/�"�h~s%L��o"��_JZ��wZ�����J��0���qF�Fg]a�ђb�h�EF+� Hd��"�ْ��W\]/���$�V�3@����}��H$��n�	UeYN��I6�3�����Y	�js)����"y3-!9��&%�e���'�q�D�'ܽ��G%K��/��֩�G�}{��[�4�&�%ڄJ��RA}�(�f��z�O��[��5ދ��O�匹�{؍����2n�'�,��*�o!��:86Ql�,L��� M6��r��Oh��s�ݹ���sJ@�'6���ip��S�Q���Eh.�3�>UŠ�5dx�j���m�^��^kT�]�lm���{]c�=3���d�5��xߟ:5ڢ������ ��!�ߢ�B��-3_�	`N���_����d~p~Uܜi�̸˓x�\3��rn/�vyA�s��B��\��d���.J\()��!o������	�Ōg�g���u��z"���.N����M9�A���M����RX�Q��ԪN�1�:�o���7i�>kSn�	(��'�������������}�������r��H;��0f�!˞Cd1 �?���� �c��B2��
t��"J4WZ)�O{�ҏt���ܪ���kv������
I�6�]q8�>"�6},��go~��� �e܃��5�tF��k�f���U5�|�)������dO�����%�;g���A�]#a�J��:��)�LU��U`�L���P��S຅���~kQ�[�)��ڍ8{���I��'�23���l�D�����*�������G�x��P	������7�J"��H�,z��s"����I��M"�ۖ%�%�Lu�O+�
x7���:pl��U�֒�yֹ�}�0s�rR逭P���[h����6_��2ێ�?ڳ��zH3`�w�_621��*���f7�.4���i���ڡ��rs�����[��6�e����O~ĕw�$D�ɩthb���*�L}M�7�/�������6[�ت�xJ���V�C\�>�1�1)�ĝ����5�����wl�f�
;�%�署����
���%�=u�^M}��� Y��i-7%����e]�fWD�;��<G�T� t\�O����d�0�����9��A=�
�F��|~��;�Rg���&8'��aу�<���-���[i�,�t�~y� ����s��?�U��mr��e�ԩ"�{ES���Ν�O����������I�WP��R�9��TPnΦ���i�&�]4k�ݗO�NՁe*�j�#��&Hգ���k9��vo<X�p�t["w�=��L�e�m�G9"�Nr��K��eA߸V�b���V�����\�s��j�ǚ��5;�g2Z�[KE��5V�=��WHxHi�Y�*�'"�����&ai*)kT�ԙ���N����֩��r����Z�9;�J�k+<[�@���?&n��)��sgǘ�~ybb�ⓑ��w3���6����q�Rr�a���:U��)�N�� �������@sd�x���(�/N�кǾ�{�������M2_ｈWR���b�ɉ۳*;ǂ|N�7�,��Ζ��u6Ć��L�D�j�1PՑ��,]��gUIhI�b���؁�	4�/����\F��������@��o�آ�� ���7�~F�!��4q���?2�΅;Q#w�$u�y�faѫ�s��NX6	5�c2@��x��#躸��[\�P��F�������_������3��A�)4������_�(�~:N���ט0u��.+� ��P^j����\%��e�Ҁ�#�Q"�ѣOѢ|N�[m*�R���G4ɰC:���~Lug⹎�y3��Lq�%!Pe<�1�b�>G�݊���Y�⨛�� eN�(s8��?�lYn�a�H�ڮ΀���k�7]R�e��G���޵�R�N���vx���l���l��Z��U���&l�F"A���L�H*R�I���#��Eb�S_;R~�{�5j{���7A�;��PU���$���0���iq�.B�՗�?��l��c�LTX����������k�a�x� ��^��c?�:徟��M$��@�rwP��/��W3���/p
�LN�����}��B�,��/�S�x�W�Fu�k��f_�˙;	ԯ�n��� ��؇}dx@��I�"~Q�����ow۪�# PM[uU���������/�R�Y�t��0����ӑ6�,�B��o[[C�̶|��B�XZR�R�Cny*�w��-��v� Y@,z�'��R�Qav>���>��]��"�v84�����f��<�;ƠrZy��
P����2,���[�_��Ͷ��q$,`$��XS�ri�C�+}q ��!�0�VR�>gʸX�_B˪��ւ��6�}�g[���L]E�i�"��Ó&X�Tg� oHXiG���z�sl��A�>%J�6�����Re�.��Cܢ�j@N�$��)��<ސ�}(����"��uH$D2��}��lӤ*W�к!�)r�T���V�a
�;Z���D�i��(G2���X0(�"
8���l�{$�x.�F'�;%@��q��Zw�����QQ�L��ve�8I_��ѯ���x��^ҽ�͍����uR����֦ /&���]ް�F��.�
4��3ǈ�5�s�tٌfWm�&�T�E3:[�t�$����$�������E��8��'��F����Oٔ6*�i�ZLS꾻:���*�-��1Hi���������8��V<ogL�>ї��g��X��AIj����^���.� A*I��Ǳ�ڶ�f�_"���8���-.^b��[<@m��(Zx���󵈑#֭�Âp���ľr�e'��'�Z"�u�JZw�T�a�f@�#L��K$��},��������N�oC��$�6����Wy|� ��A��z_ھ5�c*~D-��uUfN�!y^|��'���l4s��8�F�s� ��J�5!m�k���YK��p;k[�N	%��EL���1�
U�`�CDwY�������JNs}I��6�]�TΞ�2���d�[<;�`��(�(��� 4'󧞚<_si��.	�L��B��*n����*�1����C+��ީ)� ���:����~'�'�á����$��4�ò 
�[��u�p��3�P!|��1:7~�!x�ܙ^��6sc�7�a@q����'~{2`���XI�Gsa;m�ib��,TΓ�0��<KE���$)��*����B ��˦&��W��Gڇ��<k��v�B�S1��uI�8�o�MIRt=���(�a|�q8Y�ȴ���G�ۜ���*m�8=-�h���2�@��"�Y�}��I<oSs���N��]��eK�o~d���L_���I聜YYܻFD���[��r<%ӌ���Ԯ�<{�0=���t��R(n>})��g����q�T/<�F{\-��#F��X�!�����N[iZ��՞�k�7�b�K��?i�n�þ� ��l%4��J�-Q[�}��7UH�9�аi��nӘ��t���EV�b��%#�R̷K6�V��}q|���RZ�Y;�ͦ!��`l�����Z�P3\��LBi0o�}D�3��N(����׋����XK�3�*e �Q-U�Ց�CRG�V��Z1���ߤ�M��o��'��L@�K��AFjHbإ�y󅍍��������DqH������t��La� 5��w���n��}�L�K���j�VJ~�:ϣ7���>�T
ㄳ�Hzi�׭�${a�=>����b�`���qAӧq��G�e�5FŌ���i��is��d�&.o�&^Q����{�����y��w�ϑ�Q{�����}�P�JN��1[	ao�K�gR.���\�����w�^�)8����pT-h��8V-V���L?r�ۆ}�P'c��D2A���)�4(&&��o�AG7J�.˽��RSϙU�(�R��/b?��	��af��Vr��ϟ;_}�%�_t�
�Z"�U(�~�Th4��}�{�[ZxU���L�~p�z���j����͞i�܍�)ˤ��FMe����N��P�����5�T f�a}}�`���N��O翿h'��w�Kߚ�ևF������)$��?�m��o��L��`��=|�bj�����<m�;�JN{A���ٖ�у%�@P܃�E'��9���EZ���z��z�q���k
z��}I j��F�x�k�F���U��=��
;Z�/m�v��<�gb�I#]m�ۉA׮�]N�ѹ�)�L�M�����*��>�So�6�)/d��r���ܞ�����tDt�o�G��*l̰2���v��<b���a)��%#��t��y+�_�$��R�kW?{��Iz'���EOy��"�kR���AK
�o�}^>�X{|����ms�}�fT]f��۟��ҟpa�#��7`������ _8�Cgȏ��쟦`j$e�Z�"��al�k'zj��] hu�;"� 1ڶ'��G�MB ��:=�-�$gnW����^J_�5�Ӕ{�\��̪����H Pg��R�	�Fh}�)蛛���_��xEA���b����Sˋ��x�P���KU,��]�KqY#[�߿w��o��q���5���π+QꙧŲA��px���j>�%,�@D �h`�؝�zjA1��m1�:+z��J=m��@B��d%I��W���>#I���<��)�Ư���HhtZ;����d.Z�F�P��̚56B�|13�֋��fԤ�ۍI]�l揗B���!����HF&��l��Ƒ����Y�	�:�y��p��%���hu�a�ŭ���=���qL�6��ܿv|�a1T|! ����9m+���|���l��Z2r�^WN��G�CF�qf���D���N���˒�����[�Òq���a�	|s�Z �=)�$��M	3��s�w������KSP��y�����	T�?n�������aeD�=�� ˧�^��uAf�iO�_Y/t�jrm��l=���e.������Gr��+���[�J��5S�=��@�w��Tz����Է��)?}5��>Kds�?�ٽOD'R�������!:dcw���Zx)rU\���tD�_2+9=W��Z:�Ӵ_�	�v���E� �ޝt�No6�+�׉����oC?���֒���vT�x���O�u�����p����2�_;KϾL�R9p8���-����	�����٠���@�M`�}��7&��
�?��=�^X�y2�]��gR̹|��j����,�A}��� ~�[m��)�*!����|�niO��N�Z{h�]�3+�V�SIW�lB�������U0v�~�,)(qS�FmB&?�%��A��'�F�.�w��!�r���su�FZ�*H�b����m���ux��K�A����qEf��9���\D�����O~��-��J���P=ENz�(|R���$��N�.\���叽��h�3��D�#*&xK�g!$/Շ����� i�D S��L	`M936/?$�ޜ7�(,	�����V��֭4�te?c�H�m��}Pܞp��G�$�V#l�s�E�!n���*�eRD����m�8�-S�$D,��ύ`�K��;x��p0�;��'J��M/�h3ȵ�9�&L�l���~]���'�3%���8�m{'�d�H�
��F�T�
�Ș��F�B���la��6��uY+"�o;������1yy����ޝ��t��i� )!�͡T(1��{��zɲv�n�/��;��t��|�)9\i��/&u(tX���$�ux�|jw����B]��r`Y�TYc�X5��C$�����a[�����[���5��� zK�*�5M1�����sX:b�����`n�n��.�VP9��]Gxu�FN1���/��pQ��݆O�EO�s
��9�ݬ�oɋ����~o�X��8��w-HBr����L�ωȢ��ՙS�P��L=h�?��,G�F��|�f,n�&���� �}�[��}#HDa��vK
�� [l��*-><���$z*�Y\c{%�0�Ō��p&�LŒxr�n�-&�Ą�u^ ���C$G�`��Y�_�Ţ�$��^	��KY];0�� �If=��]>25����G��m7�"A{�g",Q ��n��X�������I�w��$�iB-qi��Q�;��m���d���:r:�1�������B[�5ci�*o6x8Y�t����0���E�C�D��9��!G ��tuo��y(�|i���ΒoA+�������74SnY��[h61�\�CU|��C��kS�3�5j�#����K6�&ޔ�Ȉ��9��.��aM�%�5�;����O���&�\��H�#_M�]�C]ia��$�֊EY����/�ِ?~F��c����Z����J�>n:���.n��W��0O�^�7;̂�1��}�)NHr����Ƶ���$�i�8���D�]�+�0Ϲ��l������@���!�~���R���L%�5�����M6����Ix�E0�&&8�2�hr�Q�B��P��mn��<����2�{��-���#7��D:�Q:K6���F�dT!-�U$�~E��7��[��m�~��B2��/���F`s#ڹ�YiWX���fYi8��$b�(w�x�ӝ�gky � �v���9l$�#pt�|�H���#F�0�'�ai版�>��{t>�K1T̍�o�&
i��G־��TE~h�;���J�׻{f�D�����yX4�Ɓ=���g=�J��f�O���i�:���,3ot�=�2��s��Q����	3/�η�/�Ij��s�m�����	F���1�n��I��l��mA��!���#j}�E6��&�ݪ��6���&�	�dh�<��x[��8�g���%y]���OV?.�g�� �;�_B���Y��)����Y\(�KT�ry""�;�N�h9|6l�n�l�b �Ӟ�r�1me����r�&n���5u��#����O@Y�q%��*��N�J��N��A)=�e/��z�=�zu��?�a,�{�ȁ�&�7�'�u.�q��m��Yg�ڠ;��s��j�/�>�Fn'�n_��<|ȍG�ݎ�w��ϝ^!Hk=�33���k������EW �!E�xΦ�D���g],�����dgq�����*�K!��<���RI�Dtץj�I\@�'>ܨz��VԎE�]��Fdf��%�'?r�d�v�W��~'#M�����^'�u��q9���e�t�d�'�wwi �%lL{ߡF�x�����B��I9+��h8�����E8�3��X���p����@"}�XM5|k�{5�"��Er���ҏ��Ȭ_����Y�%��k�[��ә�l CںgS�aż��G�I��g��N��|��O��~�M'8R?:7s�-�'��Q�By�p.�럪���M����+�&�mƳ,9�\�V�6�Qc��z屯�vx��u��\�{�)f�^����*-��f��|�4�X�.��j��tD�)�V{�=�ժc�xny	[�rr�բW�(N�;A~?�@���� ,��I��B0zQ�=v4t�\Ѣ�~��	��{	�l@��?�/��?b���`o?�UPS�F��7ѡ%�,}�W_��s����0�%�ۄ'n�G5sd/���;��ME"�W*�诐��8�@׹���s��l@up.x����w�k|׵!&�
�v9}	B�
���1;xو7�U�+�����4���眦��,�c�ԓqK��&[.'��t�'��N���^�|��x6��}��!������|��[Ky����ϟd��ČG�p�<P@(ŅJ��:���K��Q��X�iv�����B�W�nQRA���G#o{�w�bOl�t�o��DK⒛��y���k�J��i-��&*�+=����CH�H��Y���Xo�鳌;��8�WK�^�s
�d^{��q��9�0]&'*���.����w!��ߞ)������K����>�((�W&�R+Rm<rr��V��,4��hCm}1����.���?�;��Md��X�쯡 �2��?B�ʵH���
X⼻=�m��FOջ��C��^~p篬FJ�"��(��]�5��4�b�x������N������eA�����~�;@�}��te�I[�	3m 0f��er"/!�޷�Ym��Pn�A���57N���9�ù�ж�����}��5<v1T��g�5Y�ì�� �OO1zM�nfV���ڄ�OCd�� �V�	��$�X�r0s9�ڻ�`���C�A�iqwߡ?�[l��?���0�dú�?H�J�Bl=�\X�v2�J�'�8�,CM����xC��w9�6M3�w�03i�2Ѝ�n�ECbD������a�:+��O�?w�S��g����/��Tއ�\�!#ԁ�y'i����*?N��4��e�_F8G�Z���Z#ń�YgI�����{�m��-Eiݽ���8ZG��5�]-��R�������bC�뀢qJ�k���\��n�s��v��d����n���A���̩)p@r�ф��Ir�|X�v\(��\#5)K���/�r>U�)�*+�sXx ����fsM��_<��DMI��@�-�(�X[3��::����]�W����̿������.���I2���ŀ���A:EG+�%bV��Vtr�z�����Xə��Tl�RT��b���?���m��猯!%x����v��&��b��� x��`�`���t�2I�o-�3B ,��h�\�����2KI���~[��Z�02�a�;���,R�=+J����� 
�!D;����kȕީU�q�����^��\z�h�[�Vp9HeD"[g��g���q��0F�7�KJ��ֻj�	�D�v;W	֋�h�2~� ������ԑv�f>d(��qL����ΧB:�&>��ܐ#=��9��8����<�%�S����28�!�����/
�N�K ���w�UILLV��xgjW΢�H2+Ȭo��p��)����x�<�#��U���H���eYH�Wޅ#ifôK@�ʍ��~̷�
��#��S�(�@P_�pF\ý��{!���q��A����^�)m�oג�=n���3��p�7(�&]��� �'M0|���"����emkK�i�@g-T�$'y�}���@�� ��	ȮXH�3�"���Brz� AE9�uG:�ePv� �$h`�e$��\~:T�ۄ�.��&D���206[[�P���H0�o��)�{$q�L��*�FE��ۓ�T�SY�#��&�͚`��v ��;#��l��H��ڐ�eMYZ���}(e�Y�סl,bt�:v��t�:�� ���-+{��c`���e�wpp��d���n^ȱ2+��DeH�����m�U<��x���A�B�sCA��Ĺ-�v�n&}�h����l3�Ʉk5�g�^=\�ϐ�t�k�؜m�<���6iEǈ�c_F5��z�0C��{@�ƼWe��'J|�~?��R��i�B�a�ǭ�y�=��g'Zd������
g���H��c�;�&�/Pm>�EG,�{�ca���u�FA`~��K��6��MB�����D�ڇО���9���+[�$�e5�#�������!�BbK������E�@�����0n,f�������.:5#7~�\��Ƹ��W��þѰCU'FJ�y^�����A��[)����h"ou�m�iDuB�����ŉ�s!���y�2�40��
���Җ�˃������!L-l����@ÌX�*��M�����ʽ�ʀ�b�g����z�ZM�K�&�q�����B�	n��#�[�~v^5�0q����z:�j�N�����K+:�5.	����_�Y�(�d�Bvfb�S8^@�J��^}�P�D�T*��0	K�/ے ��حq������Ԛ�9�%�͔g�Q�q�d��j�Or�;Hm�-����d<��n����oϧtV�N����c̭3�lo�
cϜ�i�Y�LI�qW&	9R��v�<��y|�iDq�k��t.Q��p}�W_�^i��q��/�ZO�OY*�ƷZ��y���l��8�b;��E��&H�KM�[��e2i�6�Nf��G��l>wX~�:PU��ccx�1M�8�umHI�o*�*�.�Zml�a�hCw6ݬI�00W�sΈ;,�P��@"C�'x94�s[� -o~#�*s�\T�g�����kɩ:*�ҩA�lPנ��um�g.X���^�w@�r�S�R�zzP�1����:�͸��K2KQم�h�Ճ��{�{h\l������Ny��qZ�jUTnd<[\�E|~)�֟К=�����&��ec�
}��j ���g���� �㛎���W �$4�>Qbr��0�>�(�1��eڿ�:���y��Ͻ��k@ ^8����5� �XacI��q�p}�tRnr�O�A��ˆ	1l`-ɧ��^@x6{�&�V����<Apb�h�s�frrZ���9.����5���Aqĺ�+����k�v��-���@N�r��Me��8C���k�cQ�ȨH1�ܲ'2�6���L�.��:	\>rmI	f7�BFqC {i�W�ƺ؍���8��i�zs�R�^��w�`N9�},ɑb�p�ߘAy`�S8�jE]�T�p�TX<sh���i}=y��Q����C��������dC�,ʶСρ}��?h���r����:5Ae���#�>��:ۇuo� 8/�
 ��*<�AVvrvլ��|8ː���x�x�s��y���Zbh9	��BE�T'jA��,s����v>�85����ك����IHl�0O�����1��C��3��s�
��8��F��>m�j�,\6��a�2�]��1�d�������о��H&�7wq�����d�Yz��P����*<�����k�0PI��9r=3��yY1���eY�ZN���'�����5�x�#H�A6�ˈݐ����D��2�<�Z�J�V��8��.�D���c"!��%�W-��
�@/��>��ۭ)�c0X�#���+��\�F5��Ol�~�cE�=��ŐV5L�_����0�@�X@Bʠ�;�8E�K����t�aDRύ&�����9�+��0�s��	�V3�K�:�[�#�Gjo��㿼���Z��PLa|��I�B�a�n�������$.�I_��z�)���'j�2� ����2c9��-���s�z")O�7�I<n�_�$���c�$庥��p�v���\�8R�>3}�wX`�<�@~C���jw]���~*���;�����]3�$!l4y�T6���>Ǧ��*P]� �b��ǿC�=�	�����gW���a���.�Q}�:��ğ�A��Y'�x�}�v�sNҔ��X4BkUH�"71r� �,�!�
��3��R��B�	�&;����,(ߔb����?��u��8!��$(��ŨΝ��z����2��`��b5��y�-񃫄��
�\�!)d
��]���<Уq�P�VXQ~hdZ]��4��e���:0|Im�p��ʒ�
��K;lM(�'����_�x(�����~Y���*�	��5�t�a2��'��r'��-q��E�N�L�@�WY�U��Uϴ�
h�Zb��/':��Lhmw���P�g\^����;`5)�=��4��+�Ϋ6��~�5�
c�e�XV%e[ٍߧd�Pkc�6/7�(���r��p��D�K�#����l#.3��n����bY/-�{�yC
�o���@�6 ߌ���?G��䬀0)����f��}Y�z)��¹ =x_i�`J`��D�'�K���S�0��4�G%��?�f�i���C��qW���b�lꆟ�GI)�p����e*p$vrЮ�(�JBu�a0����#���tLt�Ҧ�Ee'?Λ3�� o��Lx�D�L�9�񱛔=5�uHd�\���pC$̀cs?U�"��B�p?����/Qö�QX�8׳�uT��A��ގc��(��7Ik���[���q;���}� t�*ȐF�!:�ʫ�T�/�G��jj��2�i�d�58 N��x%ܯ\��;+�7� ���^0]��i���Kv�ϵ�}��8P��K%�9�<.n���`�p[S�hѓ֊~r�c5�_�48o{b!cO.њ�}��P|�(3>>�O.����S�f�-��k����P�2�7s�l�|(.lj�h�s�����?��:������d�=��$�^�Mn�]�ͮr�=��h�7��Y2w� ��14XK�R����,e�Ig*�X<��fG;+���$���d.�D�x�t�Ge�m�H�/�X7������$�G>D芸�$ael8�\������!2=����K�-�	)%)|!e��F���ϲ�066�%�+_ۯ�� )o�$.[�?��okҧ�% QV�7� ����� �$S\�adB����!�j�R��5��.���d����MZ��|N�s��u�r��yɼ��h�������w A�����Eۙ�����y�ה$%t<%���rDHJ���fs�"I�i��V�R���x�k
+�Q�/���S?[*��t$�
+�͏B�J�:1wY��;Bb��)���I��g�Q�c��~�CX�+*`�Ǻ���@��]�ɌE�>R��q��D/6�A�&�3$e�c� �r�M�K��O-X�����B���D����In��L-_KRyi������2��^�|@��Sb҇Ή�B2�S�蛜au��!�Kx?����Њ�Ƨe���=#��U?�W�t��"I%����uT�ه���-��V���H:��Ch���cΟW���7o�M�wǨ��)��m��-�AB25��X�8�O�����8Z�u7�K�E`p�_>f��l� �u��"To:6�KϽ���{��Kmf�!�7�|x\�WC���+��9�������Dք1o�s��h_r��[
M���ǝΉΫM�d�]���3�-�?�$�b�Ϣnҋ�"���� 3�Q���0�/�p�]	������4���s>�Gp#^s߀E��5���6�ۊMV���Aݘ?�;����;�F1�mlb�� Z�k�6�-{j�oG����p.���X�r�e��m6��O4,�T��7�-0�Wg.#5kY��
>�M���$�1dM�O�
آ�|V8�눦�33p1r�i�t�;8���z0�����!ɂ��M�GJ�èl}����J�=���:�ڪl�p��^���B����$l�i��=uױ(
�$�򬋞�j�.L���&
�ߒ�T��Gx�|1E��T!!Xqe���&�K�Rc�{��(&r���Rv�`J!�5���蜵)c����\��%����?]/R�CM��px��)L0YW��yQ����P��ZG���<�dsB����Q'��Ԁ��� ���x*V��B�$s#�N!:;�	�e���2�M�<��z�����HP�	�`��m-+�CiD�۔Pe���c0���+�,��3VpK�+�«{�-]�9_L��k�q��0^"k+���-��N�Ŭ�C|*�R��
~���̍5jù���/��26�f'Ԥ�X6,Q�>��wyU0�����:����7�Q�����BĢ66���.V��?�DЊ���#$ �3~�?��%V���M�E��x)��L�aۇF����q��3��:���8.e#<�l3c�����"��7�嬑�F`P�8p�`�x�w�-���T��<,�Iz�R:wj1g�;ɬK�+�$`�!;`Hu�|b�,�,���Ȝ�ں	ȫ�L������ۅ��F�����.�aO��j�zn
F��?���H�[������,�Z���$8rS:�+���Hj+�y�.�y�
�M�,��!2�?�bA����M�C=X\y䉾/�v}z��d �{QM��;c�w�I�q�!d�%�c.?�<_Q_����m\��mq�mI�,V���c�������@w?o��a�7��IS�qV��g[���T̿n��[m2q
����M�I�S��J`�#�匌�l��ˇx��ut9>Ox�*�^婞M���B���!N��~w�\��P�͚���QO��d��H�FC:o�M����&�d�2�x���:M�Wf9	;I�ւ�/0@���f-y�䉞%� R�ޥ�)�ݡH���LG�v��m�L�K^�%��D�=������cVC�A2: ����x��%�M��٭��ј����E��@��m$@S��*\}����45��d��P�j>�3<y�Z��s�@�M=%�&��?Y�8U+�2�$&�w*��o��	3�Z�S�G���qa��\�VA�D���Ǌ�86�G�MRv�8X�l��)�k��XT�M��S��J��ä�/�Gpz)N���N��r5�����x�[���N���������6X�I�)�� %#��j�D���~��D�(ʞg�����&����,��4��J��{�w���B���!	���:�����w���F@bR-7�}�T�ϯ�о�y�?_Z58�X�.Z5�ͷ�d����v�\��i3��9���A|��S�i�)�b�7Pu۾�n������[F���rK�q���.�{ *
)<����B�e�2���;�S%՚9�	n���W����1�<Z:;D+qH.��������p�!�0�C����V�hRC����oD�:{�C���1uU��ڈ�ARˬs��dz��Zۨ.�"d�@(v����_k�U.'9��@��k?i�Yi+�2�6�$�۝l~:;9ue5x�uM-�f�掼�/m�	0����,��#�hy\}3��o�.��)��'K�=�A��2�`%�~k��L� :��RhϠ�����Hp��Hx��9�Ռ�ۧ����|��6�b��á���LL�c��R �ݢ�j/ \�ЙėO����X!i�jٷ{*�͇���A��[.�j�_��R�j��a��Ձ^#��o�O~���-���\鍮���ޛ��ۙ��[5`R��CI�k�e�$|��L�0t�(�5k��#nO������h���.ui����QP�҂K���s��+��܊i���H�+lw`��Ii����B.�G�r��G�q��hd��}��!�D=@�s�:�u[綳�.�i)��q_�Zc��0υ.A�y��R�x�
2j낎&+�����i@��v�uay��&�ֺ_c�Qe�6>�����H���|�M09��g/�_v�^4���t�S1�8�����&N���ا��s7��J��U�tz���j$�E����ť��������}���P+ C�䙪BI�d���J|�=<c�揣�e��g[�����I!,��\~���2U�W�q�q"��4���-�jU\���8o�9�&4[ĵ:�Oz(U�+�L�0���6k�>�v�6�3��u"qE��Tn���jap9��%�y�%�ɬ�a'��/�.�]r� ��'�Z�e�G��W]��üq7��,e�y]�B�C.���>f���ɡ��( �,�c��֝$�Gl�F�s���������.�]政uZBI���r�P��x6T0s1�$�5N~���xm���D�sA}Pu/�m��Ϟ^_�[�h��]:];�7��G��սJ�ڦ���l���&nG���D�Kƚ��,�.�[�Tu6߽aGq�LGޅ5���U}鬎���{0Wb7���]{���e�7W�.U�E��)��A�C3�w-�e#U*�M��u$AxK�z�ۦc��0D��W�n�%�O;�ϐ4��з����yg��?�S�
��u�K��4D4��o�Ź��B���U�3��4��A�V&b��_��I�a� �&��h!x��q�4�G���h^�+�vm ��Y���&�GV��@ɕU����NG��(���J�rqb�.Q>�&������)'b�FwaG��~�o�2rT�`�M}�h��c�;���䈁�X}��7t��MG�- �\�,a�N�ȕ���ZD��Px��� 1��r�0�ʘV�Xk2��wF�����S;�y6b$vK� XկD(*4{���R��3�!b �+9o������CH@ ��n���҆���{\
0& 9}2���x�N��~T�aP4�"��_B��}�#{���P������;��8q9�3�j�U
���[��6�₟�h��}�ۧ2ʍ@�$s7�Uef=��p.z��WqᲛwV��c�s��&+֬5�[�˶쉼E�P`�Z*e(��r��Wx'�}iV��	_ֆf�1�wtB!*rI��*^M�}��]�d�wk�@�6�]40�TW�F�Ru�x@�@��G��?��q?�h�L���+�Ĵ�mh6NX�*�53�=���@zx��a�H,�@����Bl�l0�D~�R`�߅߉[B���=��0e��8Uv�ix��nk!W"��h}���?�q	��w�29�Z�:tb[Nټ�{�>H�q4������&�'�tuS��ɢ�� �rϠ�۪��5cQ$��^DX|9��-�9�!t��j�� 5�K҇�d��n�	���Z�������6�"c-�d�m��������?�Z������ٟaJ#�Gw����G��+���J�'9[�?�T�i��:o��(Y]9=�z�z�\H��� ��3S/��8\_h��B4/���W����+�G��!e�]����0��r��=qí�/L��̀5E�QZȊ���K�扦R�����!�=���c���.��1x$L. _p�����#p_��`��{b9OmO�2߇��k��p2"Eu�'�����v�*�e��@��.%8ɻX�ѣ�̜�����(&�ܾ/��G�D�^$RN�Ka��@�mćB�2u�r��ʛ�������J�}��X7�.K�1�y��}�g$�G(��N�Q����٫լq]�B�("�?�G8��z[UW�j���I��3^X����
6M�z����}>FwrT�jJ�3Z�Ő�U�g�.�;ꃝg�=�)WI���Z�P��L ��A�Bp�g�"�R�?���e�*��:���䒌�����ɢA������{�������yJKlb4���X��I�D���?�U.So��mnG���ݛ��ܭ�����ɣm�O/%c�rI��
���Gj����>Ǫ���Wb�Vx�)7�����XX��JYf�̭}2��ɫ���Q�g!�ro�w&x��S~c{���$��)��OxnG8��8���V�[��k�ێy��i�\�AQUX�q z���IS�P- ���F��aI���_�4�"����0�@��
LտU�����H�m.�Q[ㅳ$�)�8���L��WE���2�b�����V���Ol��=�ZY��������L�`�uEϑz�j-�Q����.S	\�鎒�e���5��=��Ȁu�p�o��]#G�mԢ���xY��g������3�`�%Q�*U�(}ڄ���P쳮�#NX�B$�8�8�G��ʙq7��ytK[��2�����O� �{�r�X���Ge��ט/z�\+V��)���f*�4x�p݊<o}��-���B�BR��KJ�� �
l���m�����JƗW1��#���	өL���?�����p5V`��Q��lp푿O4�!�!��)��4�Q�v��s�&ZyF�n;���\����$�������+?�$�XT�$!xѥG^P+�޹��(��J��.o0+�l~2�K�"�҄�ʥR$'UYԑ��3�3�P v;qO�hc|��Ɉ{:���S���%�����������`"�2�Ӵ�U%.W�[jɐ��Ur��.�9mVL?$"豽���3j�+��{�9 ��w�+�������8�REԋQц+X(Z��y1.V£G��X�k��#\�a��_�r��꣢���ĻϬ����A�Pœ�FSe���v�@��˶G��)N0�E~���O�	���@J����P���s����j�οIB�(E�Ӝ�hb��҂l���Dɗp��H:JGk�rjF`�S�ض6ӎ��c�z)Y��.o�צm�r��$%�XC�Az�}�v���;1�AT$A��Mzϓ���{q�z�u:�{��#��b���7APpI���:^�b�$s��i��-c1�.�˞��_�ZY۹Zi�;�,����.� ~�=F�$%ǁ]$�*1N�ޯ��������}C���[y�[��&�.�3���ϽOˈ��q�?N���|v
��Ƥ�4 �9�p�ƽ�O����eG�H�ß7;$���1l�tᄛ0�>yz��x3$�Z�$cS�
|��v���4�ywQ�M����d5KA��P
#g�m(�+ �N6�?#��a�qL%%�5��k@k��'ወ'l�v���#U�q�F��:�����qa������F����7c@�J� �Mz8�$+~�D�/�iVR�]��YJ���Wj��}H"c�ٞ%����'�gI���QG����|��5?$c*)��:��8�b<#��8���>j��{���sv;e]�E�Y���*ׇ�Mt��	��V(<-g}"d�N��gb���<6о�=r�H�D,=��+�y�iaJ��<w6b
����H6j�duDb\j��{��)���- �p���:3�W���p����8����@��z�4|g�|�
#��E����x>��>d��>TB���NH��&GK
��7]�K�R�኶qS���	�۠�a�+�%@d�p��M�w�R�~���z޻,��d�œ�M�E�L��v�j�^K�}��!E|��^�+q�CLɸL|w�,�u�$�O���I��)u7I}��c��/6�h�^�}A���6�k(Z�>q���Q�;L\�4'�J��(r��I�b���ӗ�pGowX���⻥d���M����HL$�o�e,�1�G��U�b�~���YW���O5��z�ZD��$�G�f�{p ���c�M���z�t����cm�Y��#O.Uϖ:�=����fh����e�#Z�m��x<+�]�jF�ݳ@]���8�[��<L�-�Ǧ�xɚu�o*�Y�B�j^�cD�g�3��(���n]����)�-��ͩ���Zb��3%�dv�l�@�nTaa�PU�OD��c�C0���tU����̶D W��"�T7�]����5�'�<:�P4���:�� �ҧ{_�S�;���uV.m]`�s
2�l>37��8���eQ��Iɨ=Z4B�r�6}C!�	E�������UW����.�5�Kolӹ��]��ޯRD&�kQx`�f`����SAib�|��Im$�J���E*���)�	��4e
�e��kE
�'�tXC�)��$�;�f�f��*��Q��j�����'7m�ۧ��'���ȡ|'(����[��������k`�Fjw�%n5�����ऍ��q��w��r��K�AE���{	[��^����QhÁ*
P���"�9w��{�FZ᪌{s�/"ݳȰa؜�T�s��D(2^v�gm��f���]6�լ|�Vp�d��5�v_=I��r�.���J{�-��; L�=>�Rk���qh+4����4��6&'�f��Q,i�i�!h�M��A���7K@������/4~ ̺S�>�{�����Z*۠�謶E|v�W�C���y�t�g�?�L����,w5��N�zs/��Z�����)�[A{����,��;�J}�����D�a��Z��]��y�N=N�h�A߾`S"���!`] S!�"���6i}��gp�2��������v ĺL��N� �iHn#�	��dR(�G $H���+<�`S¿�GWq�,Q����wlhS#P��QwM�N{��������S{qˉ�S�[`�b�}t�����Vi���J�$5�}ߡb�,�ز�h��`
I2l��_/��T���f3~\�A�;3���s���`�!Y��1چD�8)��yW%4Wa�m�$"��������,}\.~�7&�x��mw�� Ӭoy��]J��t����T�K��:�Z�[\Y�:NO~B�~4l�a���F���ݖ�oOۋ����u��ȗ�?���=h;��zB:�c�l�Ԁi�T�i�gHh�!�8r�+VZ�qn�����g�*��Թ��G;���R��B"�����[-":_��ٟ�p�	�K�nDH�x��)|oS��JMSe4Mʒ���i�a��S��p|�6&�h_���x��������{̡u�SX8��X�&d�<
A�,��F|�䨃�(�KB/Q�N׉]�u��-�8:£�Z�ݿހc	o��v�J�%"����}��RYc?���u��2k�j\��Q �D!�v�����`�S�ɜ�]�圤2*ڨ�Nxe�(�L7SD,-}���(`]�فw5z���:�&5 �g%�z)��w6�I��X��*ףh:�H��}ItC�y%g`�1���0�9~%�$b�q���B�' "+ugJ9eS�.�2�z�R(�y��Ű���vb "_o*4�+�re���,�l3�,�H�	�i�J�=f�����؊����1?����텅l픔������%8�0ʩ������_@o��`j�m����L���O����f�mL׼k@�����x6n-�zH�2j&�]��c7�E�e�]8��N�\6�u �����ӜL#�u��u�]c&�F�?3��lB��:z��
����dʆ�_��`��8�d��z@u�)0�2?����$I�D_������6�砬%졠�x[`���1�&�;�s\,D�n^Vo7���Y����i*�.��~C_2T�z����3��g�L,�w��=���B��Y9�[9�U��j������w[-Քn�řk�ï;ʋ��է�����W�x���UB��y[<����G`	F9` فg�li"0�Y�7��<�M%Iۇ��6Zn�:	��E�k�f1n�W(�5�l�(\<��m�V !�:'K���VO��hM��ө2�D�`71���!Z�U�mdM�5Qi�{��;����� �B|<e:��<�tV��%,UV?��}\а���(��(�b��Fdq�Z��l���kmV'e��N2�� \iG	=V緔�����N�K3���^'t��] -{�1�i�	���������iCE^����>;�w�H����oI�����٧TD���r�w���e%m�O�$(f�e	o���ЁN��6Hei`�=-�t��s��o&��7������T)��	��"K)���-��7� m�����r� �|�Ю~�2����f<���T>�oO?-��v����^���4ӳ��eO-ާ�� 8U.��ΈT�8�
*v�,�Ǒ����i�V�e�^<���tsjd���F�Z-R7�d^@v��r�� C����LsT02�d�x �c;�6q�.�V|z�
������r\�.u�X�(;0��I���Ra���GދIː����i��� ���gdOŒC:�-����Q��k�T
�e]�6�<6	��,eu$.H:<�BJ�\YPw��߾%s-07��T�R(��0D���*�����P�&*mSVp_�Vq�ew�;�(+g��K NsO]P����cL�,K�S��#�|
���>�F���f}*-$�J�%�1��~Kݡ�vҺ���B��[!������Tc9���M��z˂g�[J�O�:�^�N�����Đi��ce��$��ri��:�}D7���F�@��4�Vw��T�S�6�=*h&��W �����[�Y�.ʒ�5",C��qƾKeH��q��?����W�^M-t�m͊1ڡ���к7�Ԉ�0[���J��`,R_�co
X�T�^Svǲ�w��EZ��V��*��χ8�Q,<��Bd�yRB���s����Ï?�w� ��s����zcJ�Lk���?R������1ߋ�let����.�m�A�/�l(��iޢL�y8HǬ/̢����yOC�99�,l�P:����X����W�5��QS3��z����9�@��S��Gh�,���@�X{�{DH�(��H��=ٕU3!����j��!�-'�Z?ja8?
�no���j�)��ۍ2<�Uw���ʆҴ{�?x1��$x�����f�ȍV���3�8`z���9ŠáUB���y���ջj�(���)�Ʉ�Z#�����\��R�FP�Ε{p�l�C ��!�~�
�#v,�����Q��^Y����9X��US�tҜf�i"��[�r��(��3[��a&�mH�N���ɹ�[�e���>_}�ۙ�N!K���s�Q_�g�rrm1R�Q��`Vv����Y�(V���n��1�5��I8� X]�ۈ�y/7�x�lQ�z%B�X50��$�h��覥�50����=i��|M0�ۂ,c��a�Dx�#($�P�}v%ג&�j\om�|`-������AD5�"-��J|��rȺH�d���i�V�zv|P�߰�a۲9���x�'�Pu]E� ��y�O ����EP�j,uk���t F(�~�%oun���0ɮ����F:��1����L:�N�Y�5��Ch
)�����+BN��s��#n���C6�]�ى.��H��T���$�xLpG�i����?����'_��l���ɮC��G���-F�����шe[��nW�D1�2|�:(�*hԅ�ӌЖLN�C�b$x��U�D��*0��-�7�[q����?Ca�%���lg�����t��{�H6f
U���(V�WrQL���v�;)��c�T����gv�	��y,����� �|��Q��;RB��Ft�z����B�zp�ޗxퟩM#����f�HQ�V��=�&��_����+Y�8Ռ�]�Q�Z�z��gS����IF�����YJ�`�f|�q�ܿ���k+�f���r��z�H�����h����JckQi�*�H�IL>D���k_�i��,��J�P���N8A��0.:B��K�
�S�����9�(�i}�S��5��C�H�.a�&q�=�)�^䗜��}�J
�˝���Ň���+��g��������)U�x�t��T���E-t�8����b)O�0��ޟ�$�P(.��a-���҇��F���A�%�q�)�!�2A��!�ZA�+hU�f��T=]e ��%�o���s�,�E��d �G���w���7��AW�<�8{��L���\d��7<���i_Ȉ�%�<X�JOԨ#4���u��(��M}5�fhF�� 8B�	bi�����mv��KӨ�"GF�q�g*�`*��3�'qO�?�L�:�l���|z��,�L}���=n �C%`��G�6�"�T|����ݝ���
�������̪���w�x=*eaS�T��y�#�q�]���R�gk��������v��$���s|��o�����<S�¢�l0����gW�&�fs'Ls.px���p���֚�f�/�AR.��Ev.y�)�-�������'M��5� �޶X�����{�������q���E�I!m3p��?�&(���2�����^vE�[#ܯ	3�z��^
�9��4���|��:�d����0�X��R��>Y|��>�9���=�����nsG�K��<��������[vͺwu�T��DI�zf�a77Ox+��U�q�W�,���w�VZ��ʏHu�r@����W�i��zĈ۬�Y��T��flnPc"���E���$9�x������A��1�`��Ӆ}.Vp�3b5�j�� (/�qv_�")m�+���;ÞÍW,+x�����,+	����M��8��s��94��_�R��|c�P\X��l�ޑZ���'���m�u�-�=Ԥ���zV!n�.R�ϜE�f�؆��~Y�%�/m�tU�:z)�y�*�8� z���"���k����O;��{�+/&@m1�A���l�����y��?�T�@�f��4�Q��!~�]Lĩk�*�c�$s�N��𷓐C�MP��su>?�&�����BYzG����0-`K�� �k��{��v��CʎQD��N���3��MȄ[��"ֿu�a�\ԃ�;��n��&�f���,�  �B��8V��������� r�6�������Jm���b�*YW���El��q�^�qB��f�_j3�wO��5���Z�%ܹ��b)l������+���W��LH���[���P��	�n���}t�W�K�5�c9DQ��������S�h�/::�I���2!]fQ{]�9&}ȳz��(s�Kl�&���$t��\��2"fT�c��O�lb*�h%�D��!o)V��)�'�0r��M�0�RmK=�1��@D�͌ܩbeU�'/A�nR��TD<�`�w�?0���q4�(N��x��b^(�덗hP� ���F�f�wg����>�s��)��;�AP/�3Z�>��@��%}f+|!&�N�w�A��K�#�2�|����k1_�Wr
cU!����Cz:k�9�����;-�|�*f�j�!;fv��˜�{�4��H��-�T�s��b�9^x��?�#�y��A�w�B,�=a�`x�����$�%66{@@�b�"�K_Q�>��yU-X��h�'��-
�����?�P�2�R��b�޼��9�e��~!�X��v�*k����B璶�]����'5�*'�5�����c5ϱPqIgo�4�h��?���P~��o&�<����:�mkl� �'�har�_�z�2o�n1v��V�xe�t��r-�h7G	�J��P<}H�ZS]O�f�
, ߉CM��͆\��%ؖ(W	(�� 6p"��,#��\k�X�90l��'#�|H����|V4��[����5�-EF��~Z�8^6C�n��\�چl�����Ȧ&�-GlT꫄����S����"�Q׬.�X��l ���38i��B���>S3�Y����s�Ӷא
�:{�
}��+�mw�F��ِ}�W[g�	�w�^��@�x6e.��M03���q�?�׌3M�.!�(>�p��s�:�1|8Z�.���o���:zU��� �&�������5]Y?�/4�E���J�.��ܨٔ �;���jE�ڞW1��s��K�G��q����7Ԇ�y��4-GH��l�/���H�7�6�q���?R��z��d�G��{��N�5�)�y��L6��8*�Z��OW�\��-~:�lQ�Jj����S��"�3+���bޗ��rS)Y�Z�h��'�"J��N���嬨��]�ȕ�4���ӳ���0�X�g�r�ԉד�*�v�q��`0t��d}���1���5~D�F���T��}�Y���b��u's�}��2D�%.�u�9įw���C?�N�g�&�c>CR��S��.5�jrX����$���U�~�>��c	�Q�*���ۗ0�oY�Y �� ��t�#@��ua�����d�b��k�}�(�����!*��$�0{T���� h��i��:^Z�ޥ�I�>��a���DϿ�|��?0��7ne��WTy֣�(��࿱�o�%T��DE�o�\W���β��ÿLѦ�P~F�3l��K4FMЉ�T������FC�`�\(mr��bxg�Gṫ&Y��� ��é�|��&!#"S�X:swM���A��t�D��'Q�@#]*p�ܓ_s��#�+y3���jP�w��R��Z9���v���X	�ה��+�\a��K���7�"ς���gr�_����������-<�n=�"V��<��79�A��ՆJ�ig�\M�S
��t]+Wu��*Xs<:
<�?tAF�T�RS�˴��#�{U�"�rˢ����7D��Y�\&�P�Z%�Q���e��E!Cε���C�]R��s�M����Z��E�hʹ&©'�Ŵ8�����O^��3�
�=��x;���"�T�y����PFF��Z�jV�C���v�*r[G8��C�~�#�X�5?c��Hԉ(�Z�0�33r�뀥�M���|�1�p��v�j�a��s�a�����������̺���������(]��e�ˋɫh�6��FV�:���jk䞾��, �t�gZx i�⸆��#��7�D�?�n@S2����M7Żʩ��,��� $9*x���7��8��~S�����N���3��N�$aܥJ�4���U�i;?P��=�W󡦞���$�|����Ñyu�u�G��d^��e۠?SUt����"�f���m��}���'Q�R����W�<?:Ou��fl������ĽCF6�l&P,����BwíXi�G��Ba=��q^ƍ!S|^����K�b{���.M����Ω{�%c��3s��O���:�$A��K"� }��Un�W�����x���-B���[N9Ю;��}�8�봯n��Ѱ��n3����!�߲\�Cۥp����@�����?hu��)X�k/��������n�Ga����6�`W�k)�4����ko���J��1.	`�sB4а���!�����2�d�II��J���N[���.����I�P���t�g3x[b����e��|
�i�K~�Z�����3	���X���RI���)GT� 0�$�¢ֺ���r�ˑ]13�#I��x��R_��Z�`������h���@��g��m9M�Zu����}�*|��c�8���֐0��p" ��9o�l�2`9�tI��s4���)L��ZI	_ܞ�1�lv��cGv�1m��O,*����rB����4~=Z�n�_��(8�\Q4����Y�Ӄt4��L|^�����=�s�e'�3[Z@B����
2�Z��弶`f��>� �G����
�;�T��^�+��!�8`n~�l����~���R��0c-m�7�=�N��4�q����C'�d�/;1s��5��-p�u���T��	eGF��Q踞���Z��^}`��"�%C*=�)�S-�pyu�3��ⴽ���5�4T\]��,sLeBx�֕٭�q�_�<Cj�#mb;�N��$\z�����쪞~� �Ĭ,u�O��R�iP� 1�s2l�`0����umw���[=;�J�PgB5g±vD��jL�
���&Us�Yl�T�"�Wz��H`�V{����#kb��=�ef�w�4ߚ&>;HE�ki��� �3����D��R�k�	��a{�jQ�����"B����ʫr_�����Rw��E���Oj{�f�\���b1�>���3C�}��ͅe\w��|��s��3�� ��hh��ٮ4�F~nܤ~,>���ȿP�jF��0V��mJW!L5m�����R�POn��������PTO\ğ�c��S4�![��=5�۬��Kٓ�'O����?�u.Uk%I��k�u!u�~��'��S�w�֑�a��d3K
��a���1y��� ��\��n���g)��ݪ�G�8r��nS�_P�M,�*5�QjC����V������h q�ͻΠG.a�b��Ѯ4�/W̃�
,A�Ȇ��n�n��kN��T�e{��??�­6��O�I�s;}M�W]�2�4!�I -pg~�m���?�QJ07� ��g�}�Bm��dWI+��؇D�J���^�����%:'�C�r�	ǻaNE>*�(9�D!8)YzLY�q�V�U���\���Xߜ(̋�1�A#g^0Sn�+�iz�˳N���#��C��{"j��\����5P@��n]����;%$�����nޒ\���Qf�M$RF�%s��/3�Jb���x�X]!1P�ܧ	+��X[�b3���W�s<���%��
Q�6��~�� ��қ���_{��9��l�K�� ��"��.*�ܛ߸9Z�NIq܋Z��4���[976���*l�8����4���.��D���>�'�o���b��"�,	Qj����x,��&�m��[��'uL��h��f��`1�Y�f�0�:���پ�1���b�SƇOX
{�\��ߗ� �ON����B��n�w��p����� ���1sq�S�Sԍ�P(�!4I���+�"�
�$|���Ƶ�Q	؆;�2
F�N&Ɛk����X�}\ۋ���$N���ey�q�`P�X��J&��ЮF ;{TD��x�sڊr��mF4�|��A�iuޏ&@���C�~T��Z���
u�A���C�R��zM�H����� �!y��W�-]�=� ����s�	5���k#)w�c`�N�+�u[&�-�D6�Q��6�f�����|�6��߂&��D]��h�E&7ZEfTBe�i��#��cď,�7���&���}��V�,��7�<c���f�zs���\ƄE�c��= �ݮU��%�|�`(�ρ]�y��&F�RH<�����@��P�
OFP�V@8\��l��@�N��������<�Y�3	��iA�?QD"$��[�Ԍ�!�>6�SK�"G�4W�A.#�"�{@:+��{bm��	�U.&�%��XU����1�iv��͍���qH�}��q>Lz�EB����;)I�/�v灱�ds�~�ܤt'ă-��u� ͸��q�jY۱��%��.c��k!�D��E�(Vv_�s�����،��+��� b�����LK��T���:��/6���48tOƅXSD��m�ܝ��
o�C�Xc�� ��J+?�P0BB�냟:H�q�hw�ɳ)/��+�,�#V6S/J/�},�]�4��>�X�C��'Հ��k��|7J]e�#cT f�W�͓�2[��W��k<��g���; ��mZ�m�B���	a�%i��������/Ird"�eǇ��H=��H�-�j�Xx�~����ŝf2n��-�/;���l� �1�w���>�1�~��ap U����i��NU��/_�魍��8���TGW�Ɍt��B���3�r����hd(��!L��I�>g]/a�w!�Ոe�9���t#Y(,g���|!<�D�l��Q���dQ;�9cSh\��:�1�G�_]@�c<{^�5�ue,i�.��e#�a^��b�>�#�����9�޳�&5E}Ágɺ���{;�9E�����Ʋ�J��	�݇/��;u�?��c!�S��!���u�[��k���J�E���]\̠�m��3���7-:)x!7��������=*��16�ڻ��;^J�6��{0�"�z �(���1{��@�mF��F�4���`���*��?>�_�#x��^��n��t�ϩRQY��x��,<�(�m"���o�����T�	��()Ka��>Gy6ߚȰ�o�s�Mg�W�O�zi��S�_F+'`�;���������g�M�l�
i��ᖔ�'�U���y�!������� &������U�aػtzn���*�H���פ"�7�*K'�͑�	t�����]'�%�o�T'5l����)UN6��QHO~��aEo,�2�S��QDYR$CM/Bv��)�+�ͧ��m<6v4�hu���y�,�~Z�y]��Lۗ�3�d3��؈i�`y,�i�����J@��`͋�s��f�W���#���Q���A���>�18�'gc�BW��6v�sK1��}�M;ᣲ<���w3�z�d9UW�$�&?�"��؄�V|��e��H�wR��j�N��7��;d�D����[�W.J�n�����R�h��y�(����H5ʠy�t�����3��IT��� 쳤¡�T�(����0xI��%ԦT��ζH{��-DKł��$j�Wy�
��I�7�C��ċ\e'ZR�����;��k�ц��X呂y��ՆR�1ð�jl嫌^�e�7��eY$θ!��o:�.�+˯��'���a�\�F��͵GB�n��Л%���!�:�.�_7F�y�J�1���~͡Q���w���l��j��"�=D�Ѿa�!�?��Rs�/�縑�6lZh"�ޢe΀�����"��豉H�ƛ�Uz���C19�o}�n�چ�#��V�"�-���ݽU�և����2)���႖�P8쭽/��ǋ{U����<�f��ݺ" ov��gF�v8�E�*�����o��o�����Td:�Q��p����b5�����9�x���Z"*�RZ��@��v[��Z��o aBL�zy#�`��)�.Q�"��2�9�Һn8yvXV������^Bӗ�+f�Go���Kt��G����.� ��cO�:D\t�Cq�'���xR�u�.�e+�)�M�QfS���
vs���}����\>0�wNY>�p��C��!I����h8��GY�n�y�S�2\)r�HpJ}c�Z�o��Ϥ|�^�mWM�nA����$c�li|R��/�y��GO��Үzn�̓��|ᨹu�����3��l{�2u�Y��K�ʔ��b`L�G�m2&�M�vW�"���ʅou���M�-U��� ��j��x���N��&��ښ9q�ey��V{!����>'HO���}E�m�|n��^%�HM�!��p
'�{�߮�4ZQ��SϷN�ݦtq�oQ;��d�Ul�#���)����P��p�y,�:� ]�H�N�-F���@�#�ë�k�����NP�9�@�!�����`�y���+^%�������ET��A�p���r9�fA|�F	}f����*M&?r5e�P��Ǭ�CO"���{� 2o�z��j���e��|��W��Vy1e�Ήp����[�`��T3m����ߨQ��D��oY�qN�Zcl��/�h ��w��Q@��?mI�����'$?��3Bi-5[~�����e��uc䃹$^�Ul �y���!��mѯ�������am[N@��,G�ܛ��L��2���i˺�1�J(�bzlbqC�^K��]�t��T
9�����R�z�ri��J/(�Je6��j�G3[��8�к#eOUW��'A����ܶr�ʴ�Dp
�U+��!dCe�P&\��Z`��G��q��tw>)6I*lx�\g�H��ͤ�#,��I�{��ࠆ[?�xx��!c��Z�W_���V͉�F��GC��ʱY
��|�mi��FW{�D�WfşZ0s�Q�;��H�qi��*�-r~1kLj�,��7������Mh�_�4���G��v���V⣙�t����e��,eHA�*����Ą充�a�Fq��E����r�T��2� ���g���q�J~`����] Q�t ������>i���������2�g�κ�d���/* ��㡏�%�8�mp�-���єw$ �b��B:��Xn��øZ�׵���2D�[치k`�J�zBӨc/2'N�eudi#�(��Z	�F��G�h�i6M�d�)^�u�������X�*�	x�~ݱ�6��2X">lw |���N?���j(������(f���&'�̺�s4iF�^�qX@�jUy�`c �6�Pjc����@/�cjJ�&3x�y9�O_4��Y._Cq������ڹ��V.V�M�����ng#X��<ͪY9aM ��G	L��M�N-�Sض&U�y�Au>"3~�*������ĐU5�7�L�lwg���&����0�։d޼��H�e�i>)0����խ��!O:������x� H)j�C֪�7�ʇ(�'�;DP�{ߋ����ZA�o�ގ���A�*fjs� |���N�Dj�$���h�~3�1^ׂy��AL�Y��
!q\U\�Ē����i4?��&���2,�����pm�@f��1�Wn��Y�(��̔�?�䋈 �c)�w.�1*�h���sW�H��$a UE�\%�f���-i4��%��1ՉS����w-��y��>���ls��5��޼������^-��� �r�7+�M�{0>Cq�������k�t�N8yf,�a���q�=�~��HG||�X���ۼt��2�VqR_&�l������G�]J���Nr�k�i"P�K-w)r/��k稊�{V��<�\���XیK;�>	��:��0u��S��/��9�:��8k_��̽
l�1)vm\��bd�
nz�4'*T�C~~�~&�}{��&�;�	�.|��.�~k���v,�*/�/A!�6.��\ �?���&��DZ;���T�����yy�ٟ:����B�����,��tC��O�����:�Зw�؎]�u�f�\���'�$}-D66�ړ|8�7�%�{��&�+��"N7��[����GN�>�R��G�k{'����|�O �R��c�j�l��"a�s)�H�M��"��A����t�H��(���`����#H�B�!?mI�C!/e���j�d�j^L�p��/�����g�l�W��u�����_rs��{�� ����r�d�W��+4���<��8�f�)�qb_mߪ7ȸ�9[8��]S+&tJ7 u���wN�������D���F;-R[G�Y�B}�X���J��wp>���n��]��U���y���`b�Q{tCC៞�Hd��~��9�8��s\��&@�q����nXN���[ອ�F�L]�Qшi��i&w�Ó0=��܄��~��H�R
E�����V��BH6e�ڿ�6�j���_��<��WF8����%P)pwc����C�3�͚�g�?9�:�$6�����, kX�H}��!s���/�E�0��ht���?��>�*kU$�x��w}���I�~�q�*)s��,�������|�Э�w���NF�;��6���^;�yX��������]ORԅ�?6)�zb�++6�.z�����)Tϧ=d�ʉ+������&��V���G��f���� :�v;���@0��܃-0b�bE��0ˈ�-�M|�g����������TjB�R�Iч�P�U�Ě������m}��Q%e�dX����=��ɂJ[ċm�;
+<J�Y&�kU;zӣD��YD�77$~���l�t[�Vk��2\~-C����f���q1�/��=R�;?9�jm�mr������J#�]����!�dvd���(�+Cyˍ����h!���at&�u��A�I�������]��^�	�x��ĺ�Tsw��m�����*IQ�P�^�ӽ�S��A�|�\�'Z-��s�a)�eucQm=��2������`�h�����ʖ�NG�y��p����sy�~\�Dx�ws���v�<��j��5��@{����	9����8?����<�wz���7�����GKjn̡��Y�J}���_��m�U3i���\[ů��r�4[t���y�m�VX�|H��ro[���4�i�0�F��@ee��h�/ݻ*Ĕ��څ9�/�4%�x�� ��Ej>I��Ib��
�����83~7E�B9�`�AYY&�8l�'��N��a*����3�������s��2m	EXr���O������Ձt {Wb.a��VvW�M�au	������(���ؾ4u�Fdhf��[.�Xr�Ǧ��9�I�B����������ch3.�` N�"n�	��̆5���A�&~���CTm��YNA��n��}�
J��~�x�0��Df���\ܱ�
�D����-6G�Sէ2����Qʺ̎�FD�WQdC�ʯЍD��d8��("u�n,�Lz�gd�K��Z�9�2��(ܝ�� "L#�{�?�P�d��N�S���X'��
$#x��4)t���MM���S�`���;L�g+���S1-��w��h97���Y�Y㭇w0���q*���DIkv�����u��Y~�|�ԃ�����m�N�ϊN�+p2�4��3t�t��0�Qu�'�����o,A�c�����p]���kdo�RP�w�·Q��X��},U0�����"�gw� �_�45��}:)��S�d"�!�����l;\����Ȣ�{xR��>a�5IK�X6 ��@~��esbe^ç��/A���
A��+T3Y�����gl0��Ba;�~���vF���/P�
�%.��P��%�˅�����B�'H[�H�,�<�"9�薫@�Rl6}6��C��d$������
��_2�U���V��bZ7r�B��Q��5�o��w��ю��rcͺ�W@wV��q1~_(��,)GH�G���c2�Ȃ]fT���kP��/~	�O�H1�!���twc6�-70��8(�Zx�oxc�y�A}�DY�2N'���ب%�i�%�D~π��qt���V�Ⱄ�d���;�$G��ω�V`�0�.ͷ�1������ T���|b��tL���`����0TU��u���kS��w>�8qO
í�\V���l�P��w'd�_�Q�J���*2/�k.����gr�P��^��̋xW)��̟��L����7a\�qu�r�yS4�O�i"H�����+j�=�X��)^����&���U#(�:���o�v�3TI��J�|�p"��g�؛��7��n�c��2�
5"�����=VS�`	yd�Vqү�9����S6:���K>k�@���:>�0��˼d���!MP�cމb�Q��U�
,�4.z��I��:�;��t|*�5h���9�L	��
rVU����{�;�������Di���Q*�eJڡ%\z����Ep�� ��k�Ē�i��C��okR��2ߝ���IV[��K�x	�z~^|�~|x5绶2�HVx����ժ����V�L��RV�V�sC�ʵ����E]ux�A7s�t>���^��t��"�R��au)��I�	����������u�|�I^���|�h1a4����޻e66�����@�DG��/-�q�� �hT�"$�5�<�J�7ⴍ�^؜�irMa�ip�pMB��W^L�/D:#n��������?����I�kе�&���QG|��z�����ĻCŎ �ıȢg�y���*����vWs)�A�0֧��0�����X��8E���T|5:��MR/:HC�cg@@�Jg���wb�D�}�5�w��E��͇֬��KS"����j�7x)�\7r��!��a��d�����Y�dLɴ*�(o�8Gʮ!%m@/�
t��mί1x!! [&-����0�j-8��c,<�$��G�ЎwLn�,F�C����DY�M\� �����T��B�w�ȍ���ĥ��m�ۘK�f_�	�tOrm��P�%�� g��s:���C�E��{�Ғ���y�&�4L�H�Gj��.ɏg��s�����3ZZ�6t�zF#�}�WGw~��X�A����K-�E��es�DJ5(�&�����B`��aֺ��׮4t\ik��w�����a�Z:5���<�AFzn��E�Օ;fك�"���������8����� ���2rC���6��a�=K:�a�|�m�������?_/}����������ȹB�T׍nYȰ`��
V�k(�4Uz0��ͨ����O`%yr�Ś+���֓������3c�0*|gu���lt�)����-��t;z������cXG;�r�e��/spF ��hY�<�p�3���}�b�2���!��wl���\ӏ���k'�W
��)�=Wq^?#g=)������U��C��y���d��E&�h���Ղa�0���.å�0%��\��S��A��L�o��}��nI)d'Wy�N��s���3��W���\�ܴ�I�|KBg�c��ě,!��!���M�ޑ#�'Jh�p)�vLD���z��!�uAp0�as������eV	C?���
���+�9K���oy���L��؛G��:�Ҫ��V�Lw'���?����K1�u�m+������a�±*6��ŭ$�r;[�8ѓ�����S�ng�;�K���Z�$4�5�Ɣ�^Z��)H|�d:���V�;|�9���#
��������NrN?��+x���m=�}4�N�ɡK5�o�����]�Z]�lfu5y�S��B$�/δ�LA\��������r7ܗ�C�����48�8��Q5��T9��\�zm[�iQX�O�J��$*^��&*Y��CC��݅@i�(o��z�7'i_5=	�L5x}6ov���s�v&w��81ouTJ*�H,��8lV+���ݼ���������62ua��T��F�|Q�M�,?�RJ� 	?�`'X�=.�V�Rx�������(4�\��ߥS���
L0�"'��Ț{v�l�,���$W�����Aˍ�@g�{���8� y8��K˥�{���CɈ���aEx�p��yG�kN*����Y�_�k�r8���FAn�A�]Y��d����z���&���_cB\Ɵ#t��r�%ʵ�' �L־���ɟ&�V] ��:v���>O}�0�e��$�J���B�1Ҡ��ߊ3鈟�X~R��t	g�
V���3n�����彃qo>K%�_��{�=��3���Ÿ|�������q��:��oHT)��'��L
O=uK��.�Q��J�
z��wJ~5� 7w�!�^�Gy�A?l�rE��g�9XS�}�ܣV�I��!����o�� �蔒rS�B�=]W尼rm_fKү<n�8�+%��y5��V7�A~�Ŋ骸�lq����{� W�k��K��-�&�g*�o��y΍��$����I7��-����.����-U;���ՠ�wl��v�C���_i �Q�z�����=/w�y�1"-����.>�����Q4=�ƹb��b|����&ӷȧ�Ճ�9�(��2\��9t��a��\��E�۠p,�¢��Z� &�А��]���Y�g��]�uE��&�Z�wy���R�,�L2���I�����Z{Ln��X��-��U�0ƹ����������-���r���_�!�ة�O=	��ǧ6r>z�35�@`{�����^��K>��f���{56�w�-�h�|��m�4���6ȳ 4յ�KYW�	��~!9��@%���Uly�CZW��ܦ5!��C
����{w���4G�%���AZ�*Ir��{7�o=lJ0�Dv� ��Q���e񀞨�̇�1�X�Zu�b��'�F5#~��$�Q��:wQ ���5s�a�\6�h>I�=�� a��9ɳ�q��`JN�v��Ï�&?<��^E�|u�	ĝ���+i��$]�k�ޭ�(���k�t�7L��Y�N�ȕg�QkZ��2��j�׳a�|�ި�@���:�6t���A�r+`�u}�s�����A=��CU5��:p�4���&�| ��j��F��ڱـ	O�W#7�9��-�{ g�urN���������1�����w	dq*U����+Á�_�� �.��#��4i0^�@Z�� � ���U��k_���Bm!�s5	��1�'2sa>�[Ysb����>���!Jq�e�U���TL�/��~���?
oz{
�����y�����Y��h$�C6镅�z���[�=��;/*W�'�-G	��{��m\��o�SL�Ǎ��	���D.A;9T?c�9P���>���h���}[��ͨ���vG�(~� [�)�ǹ�]ڎo���uw�,�qI���[����� ���!����3�\@�����O��7��xBh�����狭�c�����sv��ӷ\�����M`����k^���[�!�o�e�c�e��ku|�@<��b�q��q���n�X�O^j���*cO.n�'��}��7l�1�C���5�1焌&z^!�϶��ث�$4-����ڙ�F�C�j�dl�E�,�����lG�b�O���JS54D�4��UQ��?��"��0�j8lH�g��_��������=w���型F��~''��PX���������I�h#ܜ���D�M�J�@�u�C���۞��9KG�T�t$�<�*�$M9S��DՋK#Zw�/`�d��Q��1��1;���R,k��
^�5$ZZF�Y�ϒ�n�\F ]o�����2y�^#�5��&���̌APT�G���5��o������6���r[����s�F�k��-�i��:3�d�a�x����4�Jz��p�����h�� ��߄��LsM��nI��?���y�7	E\"'Z�c"
F�莪�8\	]��S6vP.hGܶ�|����O<e��A3Ѕ��O��+X>�����߬|�l�,���{o��(�+*��_&o�K�`�!�7+���lr�Vԗ�� ii�}5B��u�q��_X��<��-L����K�떔:g��9��͜�3�+��/S�����|�ѵ�G���6UhQ��ĩ��!���H
��D�@�þ��n�k����hƽځ��%��.��z��m��� ��8!���\g`��o�u�x��/8��=+���{)iW�+��ʰY,{k?���i��*-�HQ(>TE�mz�u��׽:�ws.4g�YH=�Ty��=RGϋ1��g�C�cNľ�;¡�'�ɡG�!h��Z��1���^]V�^}Ͱ�����>sا:�S-��*i>Q�;* �8�����	:�^�C�!��� ��N�)�ּ�^���cu���94��E��
<@�p�R*jO0��<���ݒ����p������w�>�B��W��n?xG6�*�����p��>��7�kE��<g�tB�L���3A_���eG�+c�q�?L��^�"D�t9����<��A���R�9�2uN�)hW��n�Fpԣ�g�{���w��%c\rQ0q�G��L'�$mKCo޵#����NS����)B��"���M����$��{�U'��݋�Ik�:��C���$m�r��#!������X$���	H��Ql'8���b��,��՗c����5Q" X0�۶��t:�}���1Ә�?����u;��󉈟%a:-�YgW�W����W~0P���\��'@b{�^��}Ru�������yZحd].����k���c�I�&'�D����5�r����6a!�������<��؊�G���[�}%�6�g�^�<_<�v�ƌ1�|X[y��.d��B��r*IG��AL���=>����������t���Q�vY��q�VoG�r�.
��M��Ű��������e�B*@�g}
L��Q� �0h���~��_%~�<�
�=�%�C?Ԏ�X�Z\;8���,���o�m�x'~8?��I�6�^�������o����5�D@�!����E?�{��`ߧ
E�t����hৃ�4=�Tˠ`2�U?ܺ�bd�O�z�@��_(�ii�ŝ�С}�(�q9�s}���C��҄"�� q��ִ= ��Д^{����1��̌!��"�����N����.U��5$�.��S�v�s}c�����5sb2�L�=|~!e�E	��c0"�*8�X���W%�����hv�"�1�vA1�Xߌ���Y c��V�nD��V�}Z;g�[��ͨ��|T�Q� x-��¦Z��/��R�	�R��N �y<]�n0pR9g��'�� 3�PO>nn�:�S�]'�:��n���B��r9�M��+�&��o��BCi�Kf�<�,�|�܂o�%~!i��{�jWƢ'�T�1��hêl�p���/�4?�x$����'��� �L0}g��k;��K01]|[I���	m�t�g'��*_��mšb�	sX �!�߈�M~�n8��bۯ*o$4.ޑ��K�vE0�9��-t%��^s���S{̛,y��(�!$S_Du�2��L��V�-{�5Z0�Ē�Aw�~���H�k�0�n�g�^h�.�����Q�@a_�uw�'��7�Y�±Z(~D�A��r���k,��@ʘN0�kˊ"�F+��D
	�<�o�0��kXd"j}3޽��},��VQT��7�.�󞀻�&JJ�m_;��40�T@��E�ù���c�Z'_� \�`��_�(
/ۣ��V��
ʵ���oe ��ȯ�v#�N��O�|I���HK1�	Y��H�*;{�YJR�����&X�S�f-Ks���{�㜿\���<�|��ǹL����>4k�]4we�Z7�ߛ���X�\���l�SK�wG��
9�mmV�c|a<h�j�	�!�9�XY��\q9(B�-����P�+@���osMP���_vx���tL�w�eQ�ɬ���	���A���b���y����6E*\;ZD���[�kXO���Az���v:��A0
ƅ=�tR@���W�U~&G�p�Y���s�w�mIL{�tz����E�f'r�k��_Ng��qV2ٞq�҉7�9G�ޭ-p�t��w�Ȋ?�y-ӨQY��Ȁ���]y� ��|3 �c��p�3���V���6�o��+���%dt��L��En�S�Sw�����V�Y��%XмG>"���13���pS
�шܽ�sI�=[\��DN���5���{囹���Ө�jf�H4鯋;�Q���W8^P($f�\f�a�}2J�tJЫV�pA����
�!?Ii:ZC�S����f�V��	�x3(���k�?��F6U7��5}T��~\�φŭ>�� ����#�5?�]\{�l4�谏{a��A�+���@�l�6�Xf���"�6#�C�d��~lW�?
��ų$��n;�[�|�j7���U%�X�4r���u>���l(��JM~Z�}X�_������ESK|$gX��H�J��f��P)㚣�0�\�ᔨ���bC	jU>�iUh�-o^&���xP՚i��G.Y�[���z��?jN�_�h�.k�����ANN3�s�>�7\�+㭵,=F@�zlê�F��^��cf��w�cG?�_%��Q�f��{ա�;��ψ'K��kZe�5�@�J���1NS������%hJ��E��:7J�b�n�\�*Bk�}[D
M�^d[%~X����SP�K�e�� 8p9��q�;GGJ+��u�,������>{ �zI�t�oaB����`SvʰˮT�FH@�(1�t��Vts��:f�^4ޏ���/�fG��gdY�xش\�t�[|Vtk��<u�.��(+v��d� ��;��%ϗ���]�D�#O`q�}fw�քMá:I��f�,���H*�o�|���*uNm��f	��n,�톕� Ď���eJS��5�dUEaf����r!�uJ�)x���qf���s������'4#p�㿝]r���cq�I�*N�q�5��7�N�8�g�&��K�8�$��H@m�q�ۺ�nD��	������ }���I�JfQ�Þ��48m*4�V���/|p&{�o��#A�����i����ߔ2%Q�A�L�P����F��ٜz�5:��O�p�<b}R�+��'��HM}�<�d(�s��u���Pt�#c��eI��g���C��âm���'��_��C�*�"�����?��7ZwD�((���5������A��b?�A�R([<�]-`6�&��µ6�K�I�TH%�C3ۘp��7��m=���z�ސd�h�.��:� �ML{��9c� رf�;?��D��q�>�ǁ�'GAwn�N���ld�J̢�P�q�
l�m�AE��`Lo��_�/;t1C� !.��=��k�g͋w�����L*_Nz���Q%j���?7:T/V������Z�;rϱ�cαsm̋<NA+��a(�uC�kɇ��Y��#�����cH�kt��S\�95�|(J��G?m��pWZ�]��B�p�Ǆ\��Jn�w)@��i�n���P��ۊ��l�D� �9l��z۱�fx?�x\�l�9)^�+�3)�*{�Ly5���~ z����[`�����2��!D��V
�Kn�!ͤ�s%�x8�+��y���0(è���E�Ŗ�V�Ţ5�9���v�&�jIQ�ȋ_4x!�aV�b��mm���i������ /��^�]�>�ɵ�o��.[�4U����_B���  ��Z��~;���iT�^�V >�H������� ��*R��[���*VBY�y��T⡽l���7�5�w^Ck�X�'_��Ʋ���-��$7")e��P�_��5)X�u]ݫ(�o�"KJ���2�qo��	�A�PN���AE@�*[�q G�X;e�;2P�+�Sȁc�4o�ޝ'�V��pv-&>��4���3XuK�z����N�K�P��ݦ���!���\-����-Jڍ��9.���9^^�,囼��@�J�����#P�3��~���G������N<D�����K_��AN��[����[��n��,+��O����Q�6&o_�9I�T��tH �9�~�� K�l����l�#n�&�(�0�K[��z��	����>r��9�֡.̊��r���H���a!_�f���h��J�r�t]�ƻ�ԥV�,���<S�z�c��ϩ1'�c���Ֆ,�z�Z���z�gO��(|�-�8�_�	L1���6�k�DO؃_��?���T��Y�0�&��c�$�w�<���sb���L������X#��M+j�2����i+�U�D;��>���2cR}	���j>j�dVBw�u�-�T�y��,�ߥ�q� }��q�z�t�aj��]�
-�����PGH��_���.�)Gi�o>_8���Y�������FB�x8hg(�}E�}v~ҝ}����O�LM�w��>ԣ��!P�7�2��;��ndqY[��R+�7�d�4�I�㚱[�Z� %�l�x]I+�eԻ �;BkV���]<p��?՗�Se�\�cZ�����:(Yy��c�����K~�)5�m<���Gۮti]Rs
�������?�W%�ĭ�o����`؅�ڔ? ���d�\��Y�w%�^v_$��~3]�gQ�K�^M��3����������j���|W{�ʭ�����������JWؘ�|�&S�(ΌH7z�8vĿ��a��!�7uC�R$:�|F���*Vq!��O�|ɨR����z����˴�"�0�b�*���N��x�(H�"��Ӓ����:�3�2���Xd�ʽ�pO��wM�(?���Ʋl�I(z]P4�0�rr��W2f~ie�:Q�/	đ��Zs���������/�D�X���J��JF#�Ɨi�`��h������W�V���N���]
��	?�H���Ne�C6#OPQ���P��U�r�<�	
��f�6�b�9%���1��e�t(��r��A]�:]�lU7���.1�=85����LԪg��Bw���{3�|I,A�<�3x�+q�$�o�'ȓ-䜔�y<��9��j=	���%�汈Q���dM6u��#~v	2iHr��ȳ��V\�*��4>'��,����Jbo�<���c���;6�SgeVs�=F�d�H��u�Yj!�{��
ܘ\zS��-:?����ͫåŹz2"*{إ�[Pp����M4�7m�6�����4"3�/����>f���-�K��Ct#{>���ñ�G4�'W?��S�?㉽�~�Bmc���l���v�-7�.���ڂ��cӤ��?Q+�ӍN�G-\�NucP�����$�@�HDCh!Y���~5�qƷ��|n����O�E��H%)Z�VQ\�\��e3�
P�9�ge!��=݅���9�����fBh�����T�HH�T���2��M-��V��.S���>�
��`�,9��ޤ���P�$����m��Q8{X�'��"D�4,	��E鼡�|#9�!Zi���u�ъH9�p�
�^+w����� V�b -��?�v�B*������������^��|c��r��9�d�@.�.f�6IC��&�*�p�NI��1��,�$��IE(K������lf�#q>�Ǌk��nؔX�mc�C�vA(�4����7l7�����wĶyYN�.�F��%���qv���lR\^'Ĝ��eS1��(�(��tcf��i���9�N���_V����f��?3%�(��9����rj=[���I�յ(#���h��p��G�%(� ��@���>�d!>D�uܠ,<n�(�n
f�iR��JgfW�����(ԩ{�$�3) �[jZ
��/(>t����۩�{����2�Jvv�&�?ߞ�Ճ����=N���S�7h���H���l��z�|��1��e�!@n�Y�OY����%��U�iD�
��AJ�ܸ¿#ϝ۵է�e��A'����;�H�Y��p⧿��x�/J� iG�J�j���~�� )d���2֝�;���d�o{�]/�Bzf};����1�3���}%W��&~��{�g�!�G��=�diNX�Q5�dQ#�@�ͰR����}�+
hJ���ar��#9#�O��?$B������-�G�{ny�f%d���������c�mײ�ew����C�^���0��?J���{�˺'�(N����e?�|�()�c]��2�o��Pn�IÚ���'uڮ����W,���/������#қ��8HJƍ8����z��.�).'C�d�������(�_�7_��a����;��� �4��=%W�Pf
�Aj���oȈͳ2�oW����Q ��:�k@��U��ȏ�Aj���;�	�[�^���?�\���2��Y��N"���������1p�Ac	��5a�6Ξ?��!?��ۛ.�(��2U'��>��-G�A�l��ު�l
c�{�`�I��PX,���*i�ݭ��ݹƎ��^0����45��S-sx����9z�����1���|��&`=/}z�D�S�.���ґ�exJ����x#�g"e��&g�3b��{N����0� pa� �3��!ut0'�2���ԕ��ٚ��LLG<!H,�p��"�y��u�1��q��$��s��Sږ�@�~e��o;_�a�6�DC�x���L�4qS)�"��w�	�78"�΄�'���b}E��u�XC���f��X���K�N׍�y�?JS%�1@*a<��z�.D���%Š��{��΢W�?�X�����F�vs�'���*g��{Jf���V��/ջr��l��MY͊]�k���	���v��g=g�n�v�(4��d���ƅ H�
9r���bN�,��1ܣ��'a�f�c���r��W� �f�EI����(?L���@���gm�
)�d}/�G1��u!{j�)�H8��t3@ �t���D�������6�00_��B�ͰֱuQ�"��H�:kѧ�9Y���_�&���=� Z��q�,'��)l@�ѭH.����J�|�c~���@z�|E=?)�j�{�J���`_�t�]L�r�x��2c���"�:m9��Ǒ�zF|*��hp����ڟH8m���f���kA�O�c�X��)t���y1���wY[�<��o}���8m����=m�"�a�[�ƶ������;�Mҿ��<����ԑ�ǋp|����R�k���x�r������1�:���"��(��&z�U�K�/c�z*Ս��Ae8x���+��7�Ir������7��W���i[9�~Ȍǅ_7�8fѣ���/g=��D�=5��_{���y�8v�πWhء��Lc��D�!�Z�$.�&�j��/�c�H��wu-�L���=�q�`��@��,^ɥ�P�j����ّ����tko����g���^?ۅX�V���J�z5 *��Y~�3K�6�/����A~�*]X)�ޟy�YylK%=��B�^>M,��=� �V�U	=���h4X��:��~�a��AX���]�Rk4w�I)�<W�.�]=���Lqi�0��t��C�����W�TV3��"uЗ־PO9�|�׫���]��ݐZQ��l��+��S�Z	�e�wF��H�F'V��)9a�ݸ�	��+&�b���3��P!}G��ۭ�>؊)���˳�]N|teA8��V�ǵi�/���ۛ��-��~m��g/$�!v�W �g-�Z������ZY��8SB_���YS]D9TF�8<��8��C��t��n)fj��²�ў�wf��L��ܷ��O��=C^��I�9q5"�6%m�}&'���������(�yl*.؏ �x=(��o������(���
�ƴ���1��	9�C?�Z-�r��<��$,�vD�d.RFҥI��{���${R�
y�����m����-JjBk�N7���岯��L�;�d;�)Շ^ �Ǭ}}\-�=-c�;^,��>t]U~w		,\���s��E��2�Pa���8��1#?\�L��x��l#)� �w+Olss��K�@WJ@3�D���A��k:z�c�+iL��1mj��bp)wpK���zS�_zG.Wf��c#Y6F6B���B�nY�y�����Pԇ��ez����qL	*�����P���G1�G0��R��ӛg덛db�>�1@SЍ��s�`�j�K�Ui�d[/	g��Ǩ���	���]�D�C�����mӆ=O/ $��[oVOu�A���a&�g����~��5��tw�eL�/\�5�f������	��� ����cے<��\�\J�(�0
���Φ�7F�[$���Y���T��2(e	��R�
���Yw��<�v]�N�a"�j~�Co���#��B9�
#��,[_����ء��v@��B]��2Sq�y��E�(�%[O�m/��Z՟���./)g9^W�^,�82���t�p��jM ��:�w6��H<;�Wo}�������:*Y�%&r+�	�S~�-�x�C{8���$��`�I;��R·��8uJu#�U��O��2�3�n0�Y�����鏖3����x(㗭O=zd)|�ѤlG���o��8��<��{�L�;AS�=����B%��h)�M=v��L�-RO�@6��i{t�n�)�����Vk�s�D]�������t�������;���} ��Z�~��"��� �vB6'ڠ��N�#�?k�67@!��R�a�r�#�˽�-"�p58���9�9<s�qg�s��?���ܴ=X.l ZI{t��Ul1[cqPD?Ɲ>+�Us�܍s�X�vz޹��H⧷Ԫ'],[]xH�	���1I��P�M����+�9�`�%�&Qk8�y�i���F4r��A	�/�o3��w�aH���JM���&�v5��F���wq#Z~��x�)���.{B�����	��P��e[F v�y�a���m��A:�����*��+q�����cb��AP_̘�u�i�s]�R�X���G-�M"�E�l0�/����oT��y5#mz֨�s1�B�-o�uJR�|@�F�=>��}/.u]}T����?-�"9�;�V%�����[�6;�Au�R� �k92�f}���eO=Ч��#������DޜR6�mb�F�m}]�Q-�a�Ħ����ElI���iPf`�wX/�H��-��웭 %�Y��3�5���� �JJc��w�m�ӓ�F�Aw~��׍DgHpPvM��q2��c���\F�Β��DL�_��4�����*ݥjJ���wWd}S��ٚhM�,*g�P�od��*��m�Bo����.��t�!UU8�F����U-�x������Qd��|���{!}]ln����|��=0���NҨ>oP\K~�؄ފ�d��v�L�^�~#��6�Cߪ4۵���R������������\]���(���ሯ �ND��	C�)�:+�x���xg�;ļ�����ړ��xCt�F�2��5��3y�]�Ά(
;����ZR��I9�f�C���~�,k{v12$cǵ�C����!6�44�ߒ�4
�J)��U���{+b^F�S�~è_U8���yM��w}����W����䂽-|�ݻ�_6�ul`ef������nY�W؊cէ+0��@��gO�|;��~��)���y����m`�s���IȠ���_	z1�)N�'`/��&����<���i��K��� J޾�Q:�"D�_��J9���3�ƒ=)$}��hV&-�{��\��sa椠+��D�����;��^a�0�c���ح�s�Y�F?*��i������?ڿ�]�Л��Z(�^�`�Zv�=�7һʿY�&*�����A����]<d����ӵ�*C�#�!��F�UF�,N�ѧ�&��D&:�q��}���T�	�����I垆�6R3�繒�����(��1渠P#-��4�� a��Z���Q�r�>*#�:�O���3�Q��[��S5i82�/,h6ƈ̂�;�4�d�n%����`M\J	3��w�T��>��e�/֩s℃�L'�g�|GǱ	���&�,����GE��l��7�ڣ��~����anȵ��5F�-��:�"���~�bL��S�h�+�#�W�Ĩg{�n��p��[R_\��6�����r�?p>��IS)�!�(�2O�&"��A�
�\^"J�@��:Ƽ"���M���g��N�ۭ�W̘�	��תn@F�����y��O��eVLUUR�h�E� -�[w�F�����4�Qh ����IB�/e�>�xE�m����5d�<�F������f�l�<M�M�k�^|+A+m�s�^c`h|�3n�CZ9�ղe|3n=p'��M�*��!���%���F�
Ǫx � ��q�Ƽ.G�ڝ���u�o�V�O�^�?ᇴ�v�z�ʄ�F�l-@��?u��r��}B����;��_�n���c��qV�?�#��y�nf����֫�/����G~��^Q�&)R��\���h��(��4Ǿ2OU�FJ�"�Ž�+I�a=:C�����]TI�N�Ӛ��8��W��/����l�[�N�<Ϊ{��4�^�"��A�i>���|.#y�
h6Oک�fg�m��f���B���;�h\z!/U�;�P��(��[�D~�o�hN�w��?�.�<U\�:)��,C;G	r����yA�Ԝ�v3�mW�1�lH�%�J�A9�$�1q�g�`Uh�sqe���@�V���a�T�,D�����V�B�Sj����k07b|�Zl�R��
�8l��2G(o��r(v?.����w� �U�h�� �@��h2H�R�)<�TH�d4*.+ըzlV��yj7��E-���/�bP�{���Y��� ��]���gl���-j�U1eЌ6��H�q�����U>&� m�;����/���D1 �L��u�,�~�C�2`*����9+&�������ؗ6$�|��oܒZ��WC���A�>�x�_�����g��j$�K]��M;:$��6Ր�w�E� ������@�e��h6Pc��e`��;��]�a�b�����Һ�F��{V�#��ݓ�gjZ��6�.��p�za,��}����s^y�<?�D��u�ηחc�rW@�|��Fë�.�=_-��I��5�r�4�3���N��g�
�'�;�;��d9�t�#�4��+��n)	��m���쉥�s�.RT�� ��h>%�V�]��uX	�U4�0�kէׂ���Y���J�0N�R)v���>�2�_Yc5�Ĥ�K���c����Щ?|��Qս��'�ػ@��H?1�ލ��3����p�@0�K_�	>mĢ��z|��vf��G��j�h���
�� �/�>њ���9mТ��P��KG��V?�B�CҮa�R�z�hx@ȧ 07���=u�U
����2	LO�}*�y:HeB���5d�C���MR����;L�_��\Fڝ�2v>�,;�<�4�!bjtC�G�p$T�ز$��}�d�~S���n�}�����z*ū~eW������"^h!:�n�Fe=�R&��2S��$G o<L���ű�Z�6�d�cm��iŹ�D����)�Gg�-\�T�g8�'�TV���F�;���,(Dd]fa�9��
�����%=dn>��G�����q3`�䏞��Z=�;�{C��tQgvFx �T����&,�t�WD�Ѓ�R 2�h/Iш~C���؅I���S�Z��R"��o���tWn�%ܗ��[�t�����Y/�����j��kxd���-6���:|����l�KK°�v�G)��J͡���y�3�R��K̽ǵY��:U��F}G��AV���E�mVи�&Ms�=L�s&:��o� Z����4Ā�Ա,�� �}x���q�"x�q7���{�b��d}Ͼ�����+n�޺,҂�˯p��D��Y�Ο#?8��f��^�]du�Qȉ��+��Y(��$	��7��^^͔.\���w0��O �6�n���5��=��LI%���OnJJ�E��HS}�qZYIn0���T#�3h4�c����6C�Pui�]����.6I��%�m$�nb�~L�'���L��ߢ�}�}Uy�:v)��V��|�@�2#�~���N��;1I{�,�\��2@�(]�36y&?��i��R�Z/4�+�Z�0��=��K<�سE�q@��n���l�3-���[�|b�1N�����A���ID�Ē=2�O,����x�%�h#�?۳���E����mw�Ӑ~7�,%S�X�S��E��t�)DO�=� �f! �΅��>���ol���R! ���>n^�"���;)�gD�*�l*۠&\c1Ɂ��m#������Y"".�|>�~e\O�GPGK�����׫�QXi�/��Nt���uu�7�Q�� !�Xݠ����p%��tDI"�5���SI]8������C)x�7�j� �o�-��C��|� ���]V��,�>~x�FSY]�Xl�JL�j�E�w�@:�T�����:WHJ�dwJ?���;o׊B#!c0�H$�VR��fDE$�5��B�T�3�7�c���/%W��E���C�?�;�+�8uP��̬'�m/Hr����u�K<.9C��/˝�|�î��+8�~{���o&\�2o����X�b�Ċ�]����j|��=�GF$D�6����|j�[)Z�D��� +T�/�E�Y_���rH�=ysg�o+#�^���C��L ��S��ܗ�7���fc)y�t0����4@��c)q	��{�����U`sy�����s���Ft�pq:C��T�P�U���[_���l�9e"ފ���������Xţ�8�ȥ��J���u{�y
�b������e
T����ޫ�s�v!ъ>��7e��7+%���ݻ�=��9�z�ڙl	��q���D���,^�X�,�����(�$�`R��Z��BR�e���gU�^��K����]�b_b����l��%�%�[\��2��*�c��a�m�����ў:5��G�l r4�����:#,U��׭.��ڷ�\�A�Б�؟�����'i�*����髗����Qê3���so��x��dFc��Qxo�n�_��	?�� Ȳ%N*��7��p��>�����ܖ{7��H0�`�j)�D���Mp5��w)�v��?��%��{���k0�A ���_{��X�� Ah!�z��A�g���HA��99%�����\<����ԀT��CLX7�{4N�8���]@�ǁB��	�"��8��Dt-{!����rM��;%y�y*���S[(9S�L���Y����Bf��amg��s179Ŕ���a���Y{�"��%�P�Q{L��D/2�O���p{��������u[r�A{&$�t�8{l�w=�.�z ��)˘ϳ�z5�����3��S��q�R�8��� G��k
N�*�!�0d�5�r���*Hs��j��1��R2�6��~xMS�K���?�y��ȯl$K����/#�}�"��=וzB�0`�G� �JAZ�\��q�^:3�Nh�B��!W5���M����L��8�=�����{H`-�yRW@�>�8��|e�:���1��y=����k�rE�l)g�Y�b�Te&��I�^j�5��mgf���Ђ�aY�I��?
L�!9шPMwE��E���+P�I	Q�n&��]���>�K�B�$���T���!�䦕�l����Y���Kbk���>d+@��_����.bߞ���s�ޚ!��1������Z���G��J�N��:�m��C\]1�
u��LrF��7aN�'8(��d/�cJ�y�m|�/���&�v��uh0�-���z�g*��!�R�� u-0,�"��/a*��H$$����BY�I������#����MWqlI|n-rԮɃω,�D�U�W0��S<�le��S�FL��d�.l���ր���A��ǟ,�V�,�,$�@6_�}��&�c�����"�<T��a����`�by%�U�̔j�w�*:�n��g��Pv�G���ۨ��\�My�m���ߍ���|��r���bdD����4�!��1�p'�+��N�mG�׼�@���@�L��(��NnT�2�dH;%I1�2w��8�Y��C��@iaW�xzݺ7�4��t�ss'j� q����@���!�Z�l����,����*mF�>A���Z�nX�7$�xeрc���������+2���F#��� x�㼲��;Jۯ�̬���7}-g]>�&`�e1�T|��V�[�7��t�y'd~��`�N6�mAεa3��^�'Z�,�C����SE�C�3�v��i����G�b"Ǟ���/w����z�e4�����"�sل��\�&O������7WR�g��)�9��A��N��2M��`v��t�p.c�)�8ĩ��P�>��n��̑OFv���j{4Х��=Py��5��fs[�è:��`{1_t�+)�6�Cu�<�� �sn��F���X5��۝fX,��ݪ�U�c�!��*}�B��2�ގ���E�d8&�3ۋKNr���^�7�JN�6Wy�f4ޑ%(�;d�B�1��1b���������v��*ϦT�S�.ɩURc��)��P�c��l��{D8��N�v�9,j�6v~�oc%ΐ�&�@	�Ϫ�4�j�i�z�� Nk�~�?z�Y"&��J�T�!����m�t���8��.�0vH��}�h��	2n�'S�-n�b�5�İ8R��sz���D8�ku<�l+�%�KCR��;,�.R��~.i��X�ЂQ�D�r�)�_衐��ǜ�>�)3W�4��,T���g�����ȅ5��7���\S�/�ʕ�%ڦ*9á�;�N2$
at'��w}�uJ*$=p��7�ObJ�j��aNV� $�r3NB��|�#���A��]ݚ�~*E�3��2c]54VVx���b�ec������vxb_��1�����������O��
��L�+/}�<
�/NF��x��dl��3f)a��r=/�c��t&�.�?��=��:��Af��>�vr��j��?*d����,�ގ��)2�s|,���b��������iPJ�I�h����8�O�]V��5@�^5�܂I��?��Y���I�ͽ�G�U�S��Yp+ �\]t�E�[�������7���Å%�`yB_�\-J���<���2&'��r��A$M1�Ed��ג�<I9�
$�֎��r�j��ݏ�Ki�*��n(��9���N��8h>w�J�<2f/){k��S��-
ó@FDH���rE�d�BI��Q �J��ko뼧�t�j:Kj��"���^!���p��������0�=���z���^A'�n��K�(07��O<n����vɻ�Sp�`W3v�S}?��P ,���U�����7M���z������Ba�h����J��<�5����VF+�ȿ��I�����i����HQ�����H���D��(�]����7B��{[���3�dђd�X6U6��䄇��Y/1�&@A��ǹ�[)�
"GE]��lO�
Ѧ+���;�c�.�v��{�)�h���aO$���*�W��a�M��F��K�&��An3J�t���B���n�x=40=����І�22Q���p_z��< ���x���,ּywX�A��<L3oc�������~h_[3T��K��0���˭Si���5��W�ZQ ��!pW��h�B�'m�vE(�`!�fq�ܿG_0r��+->a�����Qp��l�Hs��EXx�ɔ���J;���0}�:t�N�Tk�9hu��		զ�n|���&X���Uձ�S�?U�3*9d���JVd='j�=W�"$�'�P��%��x�����ǈa�a�C�����'�!�L�I�x͸~HH���Q5=��}&f��L��oSN2���nC`��N܎���~�A�.qP���#��x��R�5�O{P�!Y��o}�Ў��A*y�����<������v- /�ێ�� R�.j9o׺j��t����������-��҃�җ��n�4Aw�r~���Q�/��WgG���լ�vE�F�y�e1|�.9A�����*��l���Rq���Ģ��}�00����S�)��Vˀ �� �������?�^z>�\k��O�?����J��Ň���E0fQ���	�j!����k7GS�B�[&s�2��� ^�\G=�j�
��[�����*.
ӱ�+U��-kT�w�fg	�=R�RU,�r(ź<����,�4e��6n�"��F�eg��:S��?h ���3�,b���$R�h���a�\�jy�q��E�F�A��V�|�{�K�bu� wOv>����Oc��PRU�>iJ%Y�l��;j��`R��H�z���'�&?���������!��i1f��du�av�E�}����N��o���0-��Mo/)l6@;cx2��}j+'`�|�GL�Aa��	���=[��/`F�=eįn��u/�Qo⥥�\��t��3L���J�(�����G���:�<=���$��R8�11_R��­D�ݢR�ay����֋��C�NQ��j�ID�`���G��Q�{�	��$A9}���i �`��k�Y�Έ&�ɍ�+�n���46vO��JC��:�������ӧ�S �pS�k~{{t�\��t�����)���`ʺ��F[�<��sq`j�`����W{����@إ����h0��8�;U�u���kD��0��D�"\FWB�l�].�gP�Yc��E��菘r�Ӗ~���8�9�����T�ƴ��z��d�q"����v�������ɬ�6�#�r���Җ���(Pr�i �[��M��"��QJ�xm`�IMI�]���хc��j?z�/�l�U��v�l{�hR<�w����{��-~���wP��	T��D�X�.� ��!b��6,�(��3w~����;�z3E�ҡi��n�j��x��8F��3U�R�c,�	���}t���7Kc����ٟ&#����y-C�xc4�\�MO��u2o�ȹ�Ex6Q\B.bƻZbY鴨[9�hꓜ�� y$'#̊*�&��Fώ�p�_M	B�B��lU�O#�F��P���'>+� ����٨�76����;�¸�>̣�UZ&��+�.��A𿉙���Ғ�gī���B��	�W�����C<aO�1I�\# (�%-˄Y��Kcs�_��d�țpޅl$�^�G���~��M� K��X9Щ�ۣ�Q�WKCf����UI�U��,�E2�w�*��L�[0����Y�iL̈�z���SQh^��c Qv��0�5┻�RЧK����=��]�p�R�Vr�N�u���Z��,R���5`�B���m��������2W���+��d��m�t!�=��Ҕp����޽�0{q�}	����R%���,\| \��?)�x�H����#�e��� T�<���[���?c��+lOOSu�kU��]-y䲩�3��i�%�
Xz���#zf��o�Uh��j�0JJPq0Ù+,�^Y5}lO9��|QľR^�%�A5����
�y7��W֗0f��e��P��E��U&��N�Ǣ�W�՜8 �6C�_��D�G�GXxi��C����T��#^��O�ޝD<;ƪK!-
Bj�f��r^<��_��`�@0����_i��W�U"�̲q�u�Zr"d���+�F��V' ,>C��3&Z��y�)ؾ��(O�n)�	H����5�DŢ���R�r�;�gz��䓡�\�8j�L���ιbBk��qEӮ݈B��b�6�yy�Bm* �?�lŽDp�D
��	&�r6�3-�)�����o��N!(����t��'�QR�ws2s� .fw��E���惍dЇ�/(�r�vWM.���
�7���W� ]�� ���F+eF�|����{��k4[��1L=�k���@�0�_�d$"v��	�^���� �*ŋH�*��d2��sHr񜵀��!s�cj����T�1�P��|���f%B�c�ƪ�
8��%(le7�9-���:�^q����jc��i��~�fE�����|���*�ʩ�M�b�L\��Lm{�� t�#ʌ����/N��r��]C�WW���$�CFW9�%do����[�1p+?)��()�o �t:^<��.-/*�'t˳3�5y����mF� �x�&��~� �d�v6^<�����ca��+��]7�Ɛ|e�YT�ʪE�|#��> 
-����5���V�c#t(��̨"oQ/�n4r�ņn��5~���墴��>q2��ċ��쬲��_�����b�!Ͳ��u����3�h
l�=sN:�/�7R�=2>�T����i��0��.T��>gk�P�l!}j̃(��s��I����o+���=eF]� >�:�&ޣ�`qA�0�{��?�d�:lW裙.���)�#�S��p>|eZ=
Yl恔G�u����)�w�ٳ�@�6�(#M�fBgjb�۷�Kŵ���B�]�*�ڋ`�o���̄�S��M[�jr�+�]���t�4@�=㖈twy˙�;qv�͡��p�V~)7�ߪv5�B*�RK
ϣ�����nkdP��K�M<���;T	��ӆs�x�m�u�7z�O���ӈ��L]^��52����O�\��K	����\(P��F<08sձ�ڷ��_�����\�#0_��'"n����b���} ��~(��SLQ����m�?#�+!�!W0���N~����5�:�"�ƞt�ZT8]���b�Ɉ�t��*j7�aب51Fz��}mxlH��o"G/����9�B�t�o+���|���DG	�+h-?HQ��s6	|��z���Ժ�)�x�G���J3=����y�0���O�O�q�D)>%���Dy�25fb�}����&&st�_�ٗ�0a)x����� �u8{����|(�9�����j�|��� x� _�$;���5�S���V��hzi����^�ܐ<ˇ��0�e\J�z!]��9�j�q�rH6����@��'�w��n~?�,E����{/c`�ĳ� ��Ս�!1qٌ�0��V�D�}9�:c0Q���τP�^H��~Qk����JM�9��;��걸�W@�b"�����y�{m߭�'|��q������=�Q4����r�MW���D-��*1��i��>&Ql���ҭ#b��MA��pS��Y�1D`�i�!���w�^hk��D���U�J*�$���� +������r_�=V.�>�妱��hÃ���9�������>/oφ�_�mK(A�e��~�--��ݕ� �����ޏkc�O�3`�����''p�-����h�0�C	�Y�T��5Q�j���2#�c��6�c�p^ȃ2�=^��8ɠ�$�ꚱK�������8IG�V��C�k6�b��W�݊n��$v��1 h���}\�䬇E��d;I��(��uC�'),�~����:�DƤ��p�9�)h͍CN�ˍ�7�ġZ� ��ɠ�.�RnQ��ε���Ze��s�`���4����ME�L
��L���S�r�⩚s�SX��[F��/w��0>r4d Hw!���+n�za	��3�32����q�/��	�x4!>�^{���<��f8�Z���dH��)���JM�nd��i��2�p��&T"��֐��x۬v���	�*2��/��S�d�Nc#��7IW;���4�ޚ	��Ts0��8��8��Ǟ�й���K[6)�P�c\{/�	&��
�$��M�ăXU�o�i�І�۴7@y�Clݶ_�\t|�é����Ԑ<`r��o��8��EƸb8-]EJ�Į^�243ʉg�f�%���������2�S�Z��T���I���q����Lγ!{������F�ڴ��b��P��W�V�>�q���m�y������Tj�ڭc9Y����8���}��=6�z�=4�;��ʼm���l�Ss��i0q��Bw�_E�n����!4*��!F��ҝ&��28͖��MX�^:@��2��yg4-�π	���4]��*�\�|��q}��&�ð�8�����ϝ��Ƭ��\m��h�_|��LO���7m�=��yq_�]��__�<w��4�����o���;�'`��rY�U��|q�u�M�B��>{#<��vّ�o�co���ix*�/O O䬗��1�U]���K3#.���n�ۦ}��&AJ�h�e�_���hH�Y;ٹզ�雐G����9�:�ЎDj�lAbر^�.�P]ͬ�)]R���v�'��G4�&<S�4m�a3�8>�����^2�17������Ke�43I��*�f!����C��B�9X�y������ͯ�[p�(����E_�Qg�*�_�ic�f"!�7������ �*q���T�)��5U�"�_�9�O��d	�5i��0�n��Vp]��*>+̆�s��k��i`�-��ڣ�'ˏ@r=$��Î�����$N��q�W��*�fa�ee����$#�z��k��[��z׃�~�y	�|dj�z!��m�!����P�T+L�诓����r [�h�9��pz9G's����*�t��%���@
�/u��PX�?u����5�cZ,3)�{2���>���ω�Ţ�c�U��{�h1lXD*��%��]콪x�r�H^�؋^�h�"�e$������{������q�ΗN:!C/$t�h��3�')��A��Aɨ�vn�Z`����Rᠺ���!��LCo<��ΫѶ���ݟ�pB�<�Ѕؼ�%����Ʉ�}��
�y\�3j��P�&�F�k:�&�k�S�p��s Xù�&���x�P5�'�k`ޚ偾��,��6s�G�C��NWf�<��:��0��	/%L�S2}ͳ�E���]y�KFm<S�$��mC=e��M���w���h�;���w��gt@�?7�k�)�0S�^V�]�`���,/ң�qVB�=�L����5��%>�:V��J�1��o�uh�+��p?[��F$��k���Ş�!����ع��d�x�oC7[%�����'�e�h%��4�F��+���zNT��a�}���ɶ�G|V�ɍLai1�HN�&�x4�2����Ƕ:6�����x�I���d ���|��bk��os ~9j����M��U��2Й���� ���� z�2u3�M	vTC�>�/uu\'V,���9*��w�LNHX�F�$7�7���-�_�Y�m�����w2
+�@��`nlBr�%��_�4.W��M1�?d-5��L{�!����fw�L9�+;��F�q��ї*�~�,`�	�L�۵.`��@:b��Y�]��� e4b��=�p�8���9Md��L�����ҝ�zN�"#4X�o�&s�F�~�r޶��Q�࿡��j���g`�j"�a�ʇ2�*����K�tu^�#�H<��p�	�����ˇ�zoa��J���C��0T��7���=�{CvD����8������ѡҕ�dc��v���Q�1�ێ	�%�[��z8/���J�����3��P��&W���q�Y��!���[�lE:���Y���b�J:�˯;����x�%�ԃ{�8�gl�����de�'Oћ�
��J\�7�/��;I;��5��y$	��nW��r�A�w/9�m +C�-�m�����{6]Z!ǻ�E����ye�p���`(����јD%�����L���D�Nk�h������%�(k�	� $�xd6}ۊ��a��GF����.W'AwH���c�n�)�i9��Ɍ�����j�0 �&�sr?2�zRZ���tJ3*
�jl���q��=<h�q�/�"�ʮ��*� ,�� ��K��yҙ�D�B5�j� H_�{�C&AVw³�kļc�D�M���!�>`��6�=,�(��IY�ْrR��6���=@�W$"��R���x�Ğ�m�{{�cK��#�9�6��[{�aՂ�:�n���	 d�!pԷ����hQ�������q�NpE���t��PP� _]Ƨ;o)�� f	.[_zw袥�w֛��O����S<t�����j{������{�*��#tDp���?��I��Z0tt����Fm�%�'*�27�A�
6Emn��Kp�
i.XD�9�,'e�h ��F����d����?n�.��i����f���~ n ��	�A�_-�w�7y'Zk��l=�%-�VqbZ���ȃ)r$
��q��^ �� GS�ⶨ|�fr<\�����Sх�.b��09'���%#kmʷ*���ۮa`\4��4@����C�����~E���fK�
�Զ�^�c��.��@��2��2Z�BG����+�������c������}c���}�ZM�G�p�w �&�ڲ��,o+RS������vG�ևH4K��m��X�f�&�� -A��*��m��r"��Ck�J(��H'�c|V6o�#��H!;ipNm��-[�<�Ou�����~Є9LXХ@��(fy�|X�n�ԠF�߶B��^I���)������^"C���ُ�-"dѭ@v�[Dmr�UG�h_h��T~S$�� �OB��ERL��u�.��Qea;{��jڨ��q���mͲD��?ۊ�X�m�.2�r�+�S�i��3!�3�_k{UIq%�^c���(B1vb�����C@��ϥ=x��l�N*�,&�.���N����\*Ht���Ӝ�I���!�m��Eh軞k[�����e��F6�"�>�,ŹϚ+��E�:b�y�m�1
����Q�A�%_=E�����J��]N~1�dֶ�9�8�i��͏�G��׭�3J�m,��[����c���8sM4����@���ۿ����'�gfha
�u���6vЙ��(��1��\o�H[d�j�[J�w�|/�+]�r���P���v�Pҷڗ*��b^�����m��o/|��Գ��2/�qiW�~�p?���^R%CIc�B���s��`D�m����KgCC�v&I�p�^c��ZKTќ=B]sƌ����7n.9>z7�G)"MYT�Z��zCh6sOQX��F� ����B��J��!��CW-e�&	#����9�30!ӯ~���<�l�)0���̘�H�߻�Ys�:����f�s%R��48�&z`�Bd��\c
H��n� �9S^��!h����$���^�bd����ي�-�P�]�A<2.e[!��c��&��E,���<<B�=�owP� )]��BK���6�� ����ɐ�&�õ��Q{�\"'��;�RTA9V�Dz�`u�o}�!�/4� ���.6��A��A�X%Cx��m��*CO���:}���zYf��`�r&���FYP{�#U��`���ትdM�Am�oC:	}�+�8�_*zn�$K-'Og!h]t�!�M��"��/�TK+A%Z��Me]���2=`.��?��k?�F,�.�V�\iW��%s�n�<�r���-��ú�Sq&ȳs�s^|e1� 
���;��V�g|���E��6�v"��P���!��
�Wx(x�s����.�d���Ƶ��([r_;j����Y��XBz�>�8T_�D�s�:����uMi����K{�"yNȿK,K�Ӻ��wH�z8�R�0_>��F�C��\E���X��s-�����~����������d%�u����N�S�p�WS�J[SPg �,�ߛ�i�R$k��5��Z�Cj��/��IT�Σ3Uxڶ��õ��g�v��\��vX��}����u$��_������@�*w����Uݏ��d���N�K��a�-N����ķ���E��`�����&�U�L�~��43(�O)(0e'�tJ#H3�W��<�\�Z;�="�Bے�g�2�N5ag�&�����Y����b��L7�]��]4K��2�"R �O�1u�u�H8�璱��2ʆ��5�G~`��J����Uz�¡�����:-^h7}e�����Gu�;R?�=�<�4���⒃���^K�g۵��phD|5ؿ^V���� ���`��rQ�y	PL^M#`�l�~�`_��G�G�,�\8��
�����x�2C�Q8��J*0j������U����r��#ޢ�4@MW�5o��Ƞ�0��S�Wq&���(\���Dq�/N
8���3��4Fʬ�g��Uz�/���q��β^��Lp�'B%,Os%:nm��؛��r��ZD�'gΙ���kͳ�E@�z"AC'�u�G�o�]r@@l�*69��<E�1��Y,!9�Q�^O���b\{�����O 
��rv�W)_oR�n�c����π15ݰ�E�`��VS"k�/�[3��찀Į�	G�x�{�3�6�ӜZE�c��i�Pe�����|�f`�+�+�If-�σ ~�E��x�F:�U��l�.��	���M��r	!�C����Rzg�xxY{�����7f�~��u���~��(�#�iY�B�C�h~M�������P�	��	*�?{��.<�������_9,��P���'��vVo�(�}�@��7`��~�g���"�wi96Z�Ŝ�O���,R�"�#f#C &�4�������:zE���88��`ʇ=�}���A�6�%#3BB˶�iI+x8܌��I9\����0��6;�=��"a��Pv�J]\^=�,m��lb����A*� C�g͍/'$͠�|���+��;�6L���k�oiģ ")���Gs���=���?���Xlto�j��������%i�]X�۟
Vڀ��0�7�"9�`q�J�H(N0�5QaQ�.U^�M@(_���� �����+��r�5f����k$�ѳ�ʽR=��[˹��'$!*�k>��X����Z�k�	��79�c6�+5�;8��g�T����h��\PZ:��|������Q�E�&��KE��87�ą/���X�$�߮x�:+�lp�h{ӽ��g��[?�Y�~<c� ?5�kc���Y5��$Gv�F�o���<���,�:?
�6���q)^p+.�i�/S�K���w���C=ݜu´�h�L��h�:�n��(F7]�¯�Ò�t�|��b�E�NL ��Xh���p㱎&pSA��L��f������m� 4�&����KR-i�	����H�IE�~���������8�d��<{E`�-Y���:�K�����pdL����b�n��yO��.:�+x(<k;58�������]��-ڤYD�����@7D{���$���ӆ�*�̮�ې�j�K���@?��W*?���O�d��a��\���YG�\}��cB�Ӯ��۷侄ݩ����cO�ע�H(�� ����n�YM����l�b[YQ�8�A������k�Z�FG��g-��?U�[Ӊq�ĕ'�2��c�8��!EC����,��i�|��dOп��f�%8��O-����#�=h��/�' R���%U,�Hz�mc%��r˴��_y�\��(Y���Knc��z�r-ɫ��.�[�ζݼ9rO4���c neJrZ�����|Z�ѽ�
m9j�!(�}.�[�\�+-5��pI���D�Dy�a6�T*��G:a;#�d�*,�:��˫��>o~�*�o�)û�7�4�}��ˊ��ܽ�譐�Yz���wh��I�CY�cI��V�B���l{�kq(���*�����ExS�+[�T��GP�e^]��M��^}47��lOh0מIs�n�L�ӗ�҃sE<��Q?-��fr����A�����95��<o��O��&C��a�#a,%[+�S:��iHmR�jA`� $8�{Y2�(��h�՞�)٠�k��,5��x��$�����&���+���V�I�ح*�85G-�T�x�
s�m�d9��F�)�}l��YV���s��	��qR,ðp�K�D�������0Cf痧�s�K�(����}�����Uo߻�$B�� �.�x�(�{b�GHּY+Ū.�M�p��k� \���4GީVrn.��|��g��2�T)~�"�=Q�E�6
�P.a)�u��?Ge�@���L��jOP͠��}��M�h߬Gb��xP��4O[9������	J���s��K�&B��7�z	�H�Ќ4��� �'|�Pֻ�lb�����,�~��d��e� #�9���d�|A��`��wQ���|�����������1L�y��F���ѭh�?�z�j�ɞ�ǆ�7/*�?vk��\&$���ҽg�[S��O�Ŵ"�rp֣h�ަ�����`3�� �"��L�M9z���ސ��K�:��7��:�·2��+�W LA��(\�_��������&���)>���{��"I�Ə{��j�UG��B��Po1@���@�,����E�����e8.��iV	"��uRc'i�\�j����{�KG��޽�������fݫ<W�����C�@���asi1S����f��($�/�s���]vn>�#0(=�H��f�b��%�Mʱ�����O�NJ��S��\<��:�ƛ�l��� ]����@��o}��m?��n��s[��~[��|c�Z+ ��֭A����ғyOc�	�UЛ����?�c�y�~�A�,��:p��UF� �d.�@�'����Sop�E����j�Yi���I!�C��b�����>GD.\`�b����P�)�ဌ�+=z�~
����2z�8g�Es�X�Q�)_M�č{z�>��=�`�M�C]$�]��x(����\������A�St��8�g���Y__)km��>�\<?:�h�x^�4�p��o0�D8�PA�T��S��9������:.2T�|'c��0��}R���W�Y���ߙ��;m��� `��&oכ����J�5p�$�BXѥ���aΤ��n8)[Է+�㦏,<b�Ej����;|�_ըjx9�0=�в�z=(�	JC��u.�5���d?���t�8'Z�qE*(��Y���^�#g�/�:�y�r�&##�/>��$\��3�q8")�`�-�LR��;uw(J[������h-7N�At��J�9�=b'�Bc������a��H� *cD��H�2�ye�W���r�O�
񊯶_^J[�{�d���W��?)d7����D�  �����#zv��}��� ��8cS�������"�<	4.~�V�u��L��5X�usb�Ao�Ʈ_luH�8�B<��Z��D#%���A����D��l)Bw\
?�/��~rh�q	��ut�w���b$?�9Mf-~W@[�:|xة�����И?������U}ѕd�.��Ȥ�8b�� ����W��X�)��>��Ⱥ	��5ph
��N�����K�?��[f|ͭ�x)�	2?Gpݠ�ɑ�
.*�kb7O�@���)��0;-?Fn��Ԭ�y����Z2�JM6C~h��U��+�-���ur^pg�L���̞�Ӏ��iϗ@��c��1�-�9����>b+�TІ4��>�o��de���X,l�&�������_�?r��]̌)��sWnB\	�	XeJ��W=)"1փ��η�U�%���m'�W,m���iVKV�m,XS"@Tt$ݨ|=A5,�f�k�V��ڨ;�s�}t�iv�5@VC�Q�,<DA:��zpVP�Zx$/�� ��8�1�:���Wy��m�?h_�s��%bĒ0Q�K2�7�>BGI��^�?$�h6��=���uX�;(:���u-\]�����*�s��j(i�ݞ"��kg�!� ��S����Gm��^6�gj�^
"I�,�����cF�~1�A������ӳ,\�?�5а혖wsz��?�:�i��j���*�X>뀴�B�)Ԉ$�!�e.nl���i9� �V6�x.$c"w2�V(���}I�tȎb��|�#yFy58���<(�A����~?�(m\��?��zY�-I��d��TZ�T�N����JX'�H8��2r�N�E�L��
�&��`�8@L���97����������;#橤�E5&���EN�u3��W/L^ִ�B���S`����@�����G�e��{���@Ò����О�{">�֌B���U�<��TQҪ��Ȗq��b��3����]��-o	���-�����p�KEش���5R�?��~��Q��G�";!�e�����d�=<}��u��k���(��@��K"���@��/) ���U��O(����ީ9hj
��M/��?~jF�C�`��alq�@'N��� 5��Jp���־�fq7�I9v�u!�J�}�4�cȌ�f�f�x�s �L^�m�0�j
�8��ۆ�`�&���J����*�i�� �_��L�vP5j�������*�Lx�o	#�F?��$ ��J��-S��� uW�ݙ��:�T_&�˲�zX��w.��a�R`I�At]n�R ����"r��8M��>-
��0��@�ޥ�(a���ь��x�ykh�&aU��F��A~G�m%�a��"`N�,�a�$iiw._R_N(I
n��M,��.��z��(@k��tSrIx���ܫ�)3W��7$�Ma�CVQTԒ�v�F�y��F�j$`?�Z%�@�w�ڼ�(2��)Ly��	�	��	Ѩ��i���A�M��8�sYB�vtFZj���-a,��OX�T�?=h������RIG]�0�S���a�K��ig�����8�0�L�p'5�I��0Vn��(pۆ���1���Sț�8�!�z���I"SH��Qיd��SP�y�*j�f���[``7Oj���|P�B�F��-�G�%J8N�M�ʮ�a�# ��i8��_���;��a�(ä(k� ��3�Fy�'3�Ga�9�����{�\�Z;̄�Ǌ�6��p�n�P|8d�+�'�"못������_��m#ְ�S������I~��0��ꋤ;�n���*tB+3�m�-�#��� g� �ɇ�9�$�-'�2l��"�_�z�����h����+�P�KԷȿ䩐��X8��o�5o?#�={X4Z�ƶ{`���xy,��K���^� ���4ݳ@�1�A�iba�pڗ)����~p`������g@��_C/q��ڱ����voe�59���X1b����;��J=8L�y�)º�dZ���>ٱe�i�=����K�*�(qk�si��J�)�2����$��N�".(��k|���^��I(�T��c���K'��t0���4�V�y�w ��rT�0�(�7�˭�gY��F�m�vc�������3�PS�|�W���|��N��hv����|,.V��v��q"����3��&�K����>p��`$E^��'S��wV�;�!�Ӯ1�ʞ
s׆4�lǵ��L�����B܋�yQ�J�t��2uUD���	cs��}�|����3���@y/�Q�+՛xE����&��kFm�Y��'LW����^q�筡{�X���"ԧ�r���8�!>n�<۰��͆�c"@�d^WI���/r��l�����b|��h�S��]����3Z�Uj��;HS^ٵ]��Wv��~���fB�H�E�<�\��v��΃�=yh�j~KF�8Q,�5fr�7MF�C�������R��dK� g	��Q���@����
�Ƌ*.I+t��r�!r7=y�9O4�X��)�I��A�W�sI� �̦����-(�1G�3r&%}�;cipzuR*�f�Զ�.��>�O����#n�nLDܣB(���@[ZS�GC��0h��;D�7	{�Ѯ���Y��	i��u`"�\T^ ^	�K|~Bdn�w�����
�%owu����R�{=�Q�[j�T�KME����^���a�c� f4c�	�g�r6\�p�F��6�u؎��)XvsnZ��O���u��v�?	���9��G�>m��/��!����E�m��'4�4�� B���m�'c��Q�nI�e�|c��D[�D�����5W��|�e���ǒ�z���D��.]��|aq�=�o���^Y��m�z�N���ϖoDwyȎv�w�:SW��I&%�Br�L��Z�e������ ��k�����C�F��ޒ������熛ў��5V��L��W�:�����ڄw̔3�1�'ڙ�mG�=�8?���#1a�~d�]'��<�6̯�L[J	�H��eI�� �Is͕���S��roW��z�mFIs���'-�
Y� ��c���+o\ܣM��}��!�U�eYu_��l3ꟕ���b���`��ɠ$���Έ����	ӥ��p���4f��5[�.cU��R/'ذ-F�D="��Gb�O��ŏ�;
��(H.�4��7��Z�ۥ�*�D��?82I'��c�o;�� FC��,���|@0b�Z]�g����H$f-e�a�b2����]�!2���n�E�.$o��}�P��ۤ�E���3��y�����ƛ�	�#T�&��^Ն�4���	���\n|�f��������C��o/R�Cfi�9I�}�=O~}�m\x��Ƥ��)��Fr_��q ���ץNM���e��][�m�Gz��͍�����`kEj֧*w�V"����&���R��$�
��3�������4fp��~ �������H��c~m��\n`�^5�cZ����8�n�a*�.�):�AÓ8Bͩ�v�����o�	ryC��E�C�$ NE����#Zm�u�![��/�̫�.a�B��=�)��;_������ r{/���muV���h�~��5��Q�925��^�<��"�ܐ>��t�˽0dP���)|ie�hg8k������T�m��t'���tE�q�@�ق���En}&��L�EL��8~��"6���+ ��n깥Gf�^�'P�����4vs�u��x�%,.���wC9�M��&�����͸�%���|Zj�W?�=���S���K�]��_���;��b&�6��Po;�Ǳ������������S)��eq�<6���PFi�P2�I��L�Z$
D�](�;Z3�iҊzTz�pC.w��P��8����	\Υ9`<�!�>�#%�b�3FU�u���s"�po=� ��)v2Y�d���"9�a���:d��7���?�u�Uݝ�j�[��
��lB-+�{��ˌ�_�&�N+7h�r��nw���d;}��g��]�h�@��p^ž!L�+! �"ʓ��RF����f�^�l/I�����4�p�zR�M�Sj��Q=r��Q튤�V��ڄ:�Z�f�*M��'N-��)Ă���Q�V�t��k�4�W��(�#T6!HCK��K�K�B�Ec�޲��$uO���;'�bo�-��,�TH��7����p$��C�`�t@Z\����QwWy�	]���Yd��L��?h-�S񙻹.�A�r�e���P./Z�����}�Jq*u�C����r�����Ɨ(�r�&X���;@l�Qm��e/EZU�rnSo�X'@o���nm�+I2٨Z�I
#:�9Tw�����bk�.�q^��K�@�CiQ��0D%���g�meJZY�N�q��>����Q�	ݥi�3��$b��/tم}w\�	Y9�����D6>ϧ�-�?��O�±��'"��-n�p�����G��T�^�W��RD	Y���>1w����/)�KB3�׾��J�v��X}�svG��h�8��?��{�#�ת��?'ӞJdƵT�����x$c�5�G�sw��$d��c��~�����������N����2X1�8Q2�PO<3G8�ď[ߪ������v�-����W�k�Dͮ'$E�c�Z��b<�1�)%fS���{.�x������%䌇4sv�Ge�v��&��q%5�����0i�y��$��ڸ��A/#e潫2C�Q��Ġ��OL����Yl��� �~;֘Y(�8\k��Z	�Vev0lHH��A�M9{�0"յSCͰ����~��6{����Rl��lVX�����'�5�po�@���ǹvY�k"���C;Y�2�f��uHտ�pKn�e��M�z��n���;G��	����#������)��q�x��ŭ0 ���=�߷V�b�+o|(�[�3R��&|��882�#sߍ?�B��*��0�|F豨/���yݰ��{�*�=�H��M����h��1�v��}����ud��.�1�Q���S�t��B�ݢӜ����\�vۓ��� n~'�����#b�UK1��g����IZ���Y�oқ�cu�F^�F�I��CB�;�Y��Y���-���(�@����Cy�~�κ�ff�!�b���l�� u��0]+��~���f�\|�`��t��Ĩ���C4T���!y���!Ewk���q�Z��Y�vs��M,ZH��|~����8g��3^�*�v-�^=�� O&.I��Թ��]`u�7@�TԲ�,�_A�;��@��#�O ��2���G��Y��(J��;� 	W@�l`�B����\K�\��!cw�a���["@T�]]m9���i����䢠��x��k��7��T29�r�YkG���=pT�6���&�(���p(��b��$s%�0"�su��,�t�­x�b�b�q{a|����Ga�Q?-0|�&�	u$\�X�!���l5�I{`a��em���)Dߪ��h�&�������\]�<�W#�� �_��s�#��Ӂ��Z�[�0��/�p�nu�/SU��_�� ���̗
z��ږ?� �Dvs$m$ ��>��J�Z��另��&�Z��=�����d	_��6��ڊ?B��OR��ٕ�`���ˤ������7,��e��O�P��(8�ZD3:�E�e.Dw�AIW�-}bA��(S��^|��-������|=A8LF6�)c��3�a�w)���"-+�c���0��o��z!�$���0֤�GQI���d�ݬR��3�VS�#e�`�-��W�x���.9���Vt�89,sռ>��W�7=��������[):�S1���I�j'�@d�yb�y�Q�SG�,g�𔅖�2�Ev�GY�4[\�?��<�8�t�fB����3�~(��y�l���;<r�&!�"����<��3��Ƴ%�~o @�J3~eX��
�@I��F����T�HO�q!HFQ�N��M����G�����fi�������Y� *L��m6�]3F��������k��THSSA�[�E	,�\^#�I��}���*�
�D��N��}���^�b�l��C�K�}��sgP��
�>��� 'םv�˓-��`�X��Bo�O@c��*A����2����$�u&�Ӎ޸z`���nfD�	�f�T�9���q;��$�Կ�Uy��T&j�{RQjK���5/�1WR���:�O-[z�d�x�{��|��5��֦��>���O�&j�����l�f:|V��u�P���Aߙ�oed�uώe	
3�kh�lz�Z4��{��Ǭ�d�� LԨ�Z"�u�֭��	�!D#a������#NB�aD���yy<H�)�t����
� �6�w��^t������Ǡ������n1�Ľ��m�V�,7��ǔ�8P�����cN�;�r��4n\
ø�I�����@?�y�3FfjJ)�����s\��yA�H19!:��:o�U�F�ő��6�*a�ڰQ�6���X~�w��]G���1����%���L���_U3<}O���^!����Z�p�T�M�4����-H^r������s1��xb��(��+n�o�uIt7��4g(�]��P|B0&�j�������q	3/kI	�\��qj�e��� �l4�����;^��>��i:����p_3��J[�V�W5�ua\+��ݻV5UVBD��n5��. ̾��k����w0j4 ��I25�f��j}��I��58��-�yo�p@>sq�}S5��4��wt�(�oRe�v�ڒa��Q���Ԓj�?�8�s���
eM�ɠH�a%��G|�;8g��
#�E*����u�
P��'c��uR8��~stf"Ļ�c;�6k�e[����_�T�1IY z`��Y���\�F�;�3p�=����I�Y-h���3&�涘�!޺0���>�}�&����09K�il��>�3�n��9�$�!#��/K5��o@C������2���z�y� ��d7[�Q�s ��3��ԹZJ����x/�xO����e���q��HEGMn���SDCT\,�RY_���o����; 8���3�N�)o�ks�b�����D������
$J�}��cl�Z1�$��D<�x�z�J9�&��	��+s�-&��)��)��cM�&�É��~~��bd�ԑ����~Z8�`v����R;�,�cC^��fl�7q���v��3o�d�����dm0ZSy��Ҟ��{ �B \.	��1*���8HI3�0�U5KSKnmM*4��@~?����-�#*�D�ŶRK�Z��OU�}�8��A*b���@I)D�����	+<a�:��i��Wr$3�p<#�G���q������J��Dlo���3�����T���j$���N�
>]��l���ӡf�+�xk�D*ڴ���7�p���7AnO�{Va�����H��m�R����9.V4Ġ?�_&g�@� ���Hw�C�o2����ȠE��d�%�yӅ����m�T��T�R��$�,����_ ��+��/v�Tg-h��>�꛴p(X v����1۟����%�U����Y"K��<"��H�SS��������{/�>���o������M���Uk�K	?�������QF�ѷ�!�q#h�6s%���B��C��s��܁ûW���b�����7]�)Zu�>��*��,hS�)�Fd����T'�ӕ�,H����;�H������2���W�A-Yg���ӽwT�)L^Y�
���K�4�Q�j�JZ��Tg�͔� }�A^)�|����[vƅ����I,%�wu�rr��y�b��K�!���"G��_��7w�¹�t_?��3����,�Woq�W��cA(֔9��M�wm���.M�0dâ�~�Ҵ����2e��(f.��>g����%�U:��zN�K!�%�����4T��c<���^k7WOO$���y��_T�	��ֳ�*������>����,�@��+r��9����#=,b}�K�Fo�O]��"m��@�͉ �ǘf}�/��;LR:�?�3`�=�]~]Eth>��-}�sI�I�.����2;T��V�� ����B_�����]$Z[������;}=�|ۜ�e'\W���  �g��:��yo��%�?�4�����zY˔����ϸϦQ\A�ƪ䛂�8���ti]��/;��?("�PWĻl�j�C8��Qv�
�J�ӰBffw�?�l��5f�b�8P�u�1,�<�j^3�-�t��� ք�@�z�d<������=����ȶ_�F����H���Y�@�p�Ǆk�����'@�e�*�iUB���$����\@iP�z�����r���ݑD߉����]5�;(�[h�A�k�];�H82�}=�^c��岨���My����=˖?c]�ZF2B���k`������
' �Y���Y+�<��q�?�fR���g����5[1��?�i��]�yՓ���S�gpv����m07{�[�uq=5�k���*(����G�>���U�x,l�I������j���pS�6��O�7��O>|&����RV��)~ð��70v^����ʩ?��y�S�@�"�|�Z�}0Y$�̩s�ng��jd��\(OXT��뿜��8���އ��+y�5�sT�W#�Vx(VUP��2�MuR8ﾏb<��I�p�(�}JP�D�ͨN8��x����̍*�����MI���TG�H���$�1z;R
�?�R������O.3<3"]T�*�A���&0�[��K�"�2���t�5M��!�"�]�ğD
|�f�%�������ɝHje��7 a�� �ى����7Dw�HXжt�Ռ=5kTߺ�߿8h>�c��D��bV�I�^Jj�ą�l.fTO�4 ��N�M�����6�]�t���q��*�^�}�#�>�SP��!; ,����#7���]s�� �m�C�\%r:�R�G�6{��x����eJ�6|f����t�L�U<	��di�ӚI�R�5�-�TȾTI��y|S��ߓ�.!h���>�X#���g�cx+jѼ�+e��� �%a�(\�-}����V�Q�ƹZ�Z�\j������sD
���	.�o��������c�CiP�=�K�NO!���6~7��0�h�7"�ǧ�����	��Ѯ*�έޫ�I��*/^{�+�ڔ���X��IO���nNe��>@��e[��u^u@��"L[gŊ��n��LR�1�{9l�~�+�v>U�)�㣞��"���!cB�®����`�4��o��������'��6;���U�����'Q��NNԬ I����G���ȧ��-lk1F�#��6���o��Á9�8�m�~��b,�7��>�!�_�ZI�k#=x(��7�=:Hз&�L����ϗ!�(Z-mW�vdA���Def�S�b6��_��:9�	�#�H��%�٘�R��BD���,0�
���R\����ս�Fz������0Ly;Cs�[�'�B}��&�6u�!e7n-�� ��+�g�x�P��F^Mɒ�|ZT`��\G�s>=h��/�6�\����������&9
ˢ�I�oyh�F�bX�L�ꄌ���솫�5�ԝ%�RQ�:6����?���}_�J	���;+p�a���m�Q�`�����J�@����?�~f޷á�'[ r�>�����vY��5��X,@,��uUP�8�s��y��ֲVf�t|�oJ�Y���`\�G��zSpu�����Y�f��^���H�o/4�*�ԟ���K�fw�����ĵ��+1�h�^u���M}T5�"�� 8��K�����zNg�Q}2�|]�f
�fYF��l��:�w��a�]��;ΞJghН����K�\$���Z�c��l��3|%R��FuM^�>��3e�O�F�p�gңh�F�_��K��`ЉΠ��Jp�S�1S�ꡯF�]{���w���EL�}���7ߌ���r֬�i%��R��1��j�#�@e���Ĉ�-T�-�b��5T���&XD�t|�j"2���*��4�N��}r�`��P���z�ϣ���WF��{:X-�l	1�~E���ц��í��R�k?�b�e��gg�{��yf�����}�!���ۿ���J>��e�����4Y�s���>t���[�V�lG{�njH�o��������LS�#�L�mjhL���yaݱƳ;V��m���,�-�b���2m�B9��y�,�c�|<I�� �(���`.wQ"BI��{w�jq�
��>�R��%l<����C��Zh�+�@}�݃+����	��O�)��V�(���$l1��s.���
�b��Ҙ������uT��C�49�n9���!�G�#&%���.������HL� n+0���YK�;���;�S$Iҏ�Je������@жuH�g�Ю'q���+\��c{��&��䤱�[�ܵj����2�D!�\�N����4�����y;1����|�!1C�x |k�6&��_C=�h'h�2�/�f��m)g=���s࠻m�J�Z�H%�נ���zk)��S�A]=����@�* ���m�־�[��J7��/-U�����e��6���E��+����[���^E��݂�9��FtZ 7B��+��f��Ky��fdr������ID�,�rJ`ˑ���VY��f���Germ�#/��yI�7�V��r��feVS�0bFR���"҄��q3v�P������MZ��[�V��e�䍐2	[�0䦟�}Yؽ���JJ��LEC�f�{��?2��?�q�U�������$��_��U�v����$a����.[E���`�K�Sݬ����
�z�<���W�n!/�e<����d��������y�$�� �}\����q�*)$�-Y�jA��_�`ednX]3k�{��R�Ĝ��n<�O�BU�</�֯q]Sp������ժP[Ne,/�~lUr@�l!`�W���������Y��?���qi��ھm�W�1;~�v(W!3UW<�_�)�������G�
������Z͕t�CQ	^�t�q3��x� _��.N�� Nm�"��՚���bBX����!f3%!�5}�)��$U��襏�ߩ�]n���>� *�[��,�8`٫�&�b����熥�� ^R�UQ5�3��I�2�&!5���bN�M~s<�M���#�;'5���/��ӕ���"=ET͘²���@߭p%�&���&V+���a/K\��+31T����Z8�;d9?��]a�>	b�J��ە-��B��#��~=C�r�FC�Ztݢ�+�f�N#��-OR�`��@ ͸��|������?�t��0K�$P��ю��gz�u�u[h�=�r�v�aR�>�\��K�p��g��6���E�~���)��g=��j�h&�m��-����=,�*lz���O	d�ز��lˇ�58��6�;Pᤚ���L b��ʫE�a����2lg��T�-A!��0��i��Hpz���+c�V�/Ĵd73Os��GO?-h��#ҋ"��p�=5�K�\��WS-jX�W��w6���TMs��¾,�o�$�tU@:�V�m�
*Ԥ+[������E䜾K4k���U�x
э�j�ٟ��O����E`#�D_!C.\��Y餹�A�̨U~	U���V��,q���M=B�d���v�r!��_"t�F-�>�����[T���)�G�N����H�f��e�ǧ]� �XZ�\[�C����:as���&
���S}��_cآ�������QZfQ��Jx����2�&�v$��=�:?t]~%.=5ϙW r0���ͻ�����p-'����m��� ��0&r�F/�U����2��g�v��O^.�\��Y��������.!�r�Xm��&f~��2�i��,�??����-�x;�3�O7��bg�yi��l�1j���B�u����T�(��e��Z��_��㷺��b}�Kc`������I�˞�U�>��^i~R6�%/A�\6�g[�ʫY�>~uB9�5�@s��˯O�r�G�O�����"���3�l�&���f���C�}f�'�ƣ��,/&�÷n�~�1+���D�3�Kő 4i#������Ww}�?���F"ԧō�ur��(e�#%�C���i�X��=d+�|rf��3�������ǳ�P]��nT�x�2j/˄��(�85:,-�>�٪"�L:�Xh�+�p1:Ͷ�r�j�ۣ͛!���Ȝ���,�Y+���y�n����mCYV�`�"�'�4�Mq���]�R��t�{��W�(�o�ј�/���#�%a�xn��7<I�"_&��Q�4E9|�U�PjnG��56��;�`��RxD�~�(
C�S�O�Q��I�̚��}��)%X ������ ��eh�u����I��M����D�.�
A��XHb�nM�h�=F¯���غ\a�_�U���L���~�jP��m���k��=�d���lpW.�r�΁��T��6I�Tj~���C(��8ۚ'ۗ��F�_+B���K��o�n��y0�ldH���%g0O1�~��r%��ٶ�T�]7���ɡL~t���`��I��/L9�L�k
M7��-9�®�F�������B�~w�5���/hl{��g�N������E�k�ón�(��y?�t	b8�L�6F��f`o�ǿYwo=��~��hʀ]�ҔEM�-��q�{�Q�3��(�0�Y~]�2�0�+��b�eØ!NcX�Ǔ{���	�>�\���M�Zeh?��"�r�;�n᡻_�e�
�@X�B�������ӊ���Z�?�������\�����^B�Gc��ʯV��"���@7Ѩ&eM�B����v��1��H�T:�e<�U���}:�G�ԡ�'V�����3ȝ� �^��8���a��jt��O��&YXM��«a-�y�'6gsؠXD��5?M��s��4��xq��z��`Z��Q� PM�fO�}f�2���rK	v��v���%V�9��E��-�(N�����\&co��(��썈�N�ϼwP5�O�k�Q n����t���4��cj	9H�p'5fh�����c�����?���
KkMK��g���]��%~��%���/^l]�n9�#h���"t]�S��1��f�pp"��]�<k.���T��2-z�3|�~�aY�UY��b��`c��E��K���,�nz1�̩�
���������TV$f8a,&:M�a��m�"_8�1??p}�O.l���9�^��T;uA\9��|���}�e�|2���D!��c�@;��o��cȴ~����	�2����Ki�6um�G�����ʿI����Ux�kc�j�a_���?�����w�}��h9:y@q��Q�_��%�nKG�����Ǒ�W
hB^\K^P_>�$0��r\FX
Z�:@\��T9���OQ�[�2��щ"��0h�^x�J��4����G�%j}��JwU+b�e~	DG��+�������N��Nn��9���sq�%1�⍖!Ϊѹ��T�<���o�t ���VWgv�g�%o#R�q{$X�P�����S��!��C��=��uH{l3Pwf��Af8�; �j��������O퉉�j0�{��d���vbޔ:���@H�'JhVF�h�P��yd�\��(�C9/�EX�]����39��:�Tl<��F^����#O�V.C��
^���Iǟ>��+��OR�ոw��o��ŧJ������c�w�r����pUy�ol�$���S�i2Qg��0Z�*屬��y#�g�0S�ι�t��1W�MX���fӆ��3D�k���.�K�o�3V�O��1N
wz�ցf�%�0f�M�f����ڋrMl r� ļuŸ-'g�7z�("�Q��P�۝�}�.K�J�]j(��*0��N2��E�!䖄L������<���~?�X�sJ�މs�P|���f%
%�1��膏�\�-��a�2ɿ�	5N����_3#���z�`u>����St�=���i�)H�9a�'��S|R�M�%�*�.7��)飽��W��R^J��lEƊg|��
a�eN���z7����/'Õ�v0 ���?! wO�����k	τt�.d���Ը7B�����u����O���+�XP�W���qpK��u+
��T.��=ju6l�D�$��m�AP%LΚ��]v��Nmp�#Fu��N�e��<?5#��wV��ȓ�P��{�x]�2��^�A��fu\@6.9؜��ǚ�u��"+��UO/�$�;����5��M�����(I@C[��ݘ��=b^�N����Z��F7��ǂÏ�|W�9<x�|y�gٞ΋��җ�q��z��)�_?n�vu�6��0����@j���x�m���e�i@�������!ˇ���`F]���^f��;��u�/��l�z��g���4��̸ֽ�;k���3�Ӄv&��ȩ_��0���ĸ������.���� ��x�6H۶� s]�_�VB�!�	p�}B� ���b�'���YK���qoѽ�X?�"!"[�=���-h̦�"��ө�ܓ���H_����6�eBހ�?�4sv���v��(��B����-�%�ա��΂��VK����)�nn�Wy�|75�c�M�/�Ƞ�Qe5�Q�G�GV��|�Ř߃1�jq�{��6���g��=Tpu*����D,g�+�%����{���<>�\f�{͊�F��#���Y�~�������RG+}�噘�h��
���A�W�?%����)i7��l�6��|��#޷r��@��)�[J�]�����7�$���!�L�wb����M��x��gȓ5X;dk���!7������嵅�S�,�C ���x��A�Y��������2dO%h:C��4�R�o5�j��8&G�r�n<��O�@A�G�LӚ]�(����#O4\���>4��Mn���Zl2<i���"�	s=�>��z�s����{�w)"�V�6�_���&(�U�Q�`e9������;���n�.4�&�65Bm��=;�	���DA5��5�SP���d��`�8ӂ[I�Rf��ؤy�f�%�0�f�z�
�CFX~�c������-3��Ӎ�kX��J�Ϸ�N4h��h����anh�Rw��W��C�l���fA� ������V�OߖF��ڴ�		xu�������&�쌘���_���	�Ժ O%���m��؍�	v�]� �B��A���L��eW��0A�k�˼�����lw0�3�g�{�1G��9+xM̑�Ӎ)_�����O]�k�[��;�ҀC�ya��E�}'�b����^��S�Œ�V���C�o�q7A#SH��׹��c��B�pp{�e���8�l b�T���j1&}�r�N��ލ8�9�/!4j)�,s��sY��x�h��{K">��f��đ�8��L�Ҩ�Oi���Fx���J���7����c�_]��2&X���f�b���� n*��o���B��4�q��h:�&mJ�8�SKQ6�%�� ����ܻZ�ڵ������+L���¨NO�������29B��>��l��|��%��ؘ��Co�p�u���2pV��Z(������h�]Kͅ?�*��Q+�����	uzN����lYͼƞ$�~�=��>��*p�����ޓT�r��P�C��Q�
l3��/͌$ΖY�O�5�>��y��)��,���D���=�]	(��DB4y���I�/7'�B*����Z�A�Ѣ�MK^+.:��=lK(>����
�ؗ�ܾ��4��{A��4�}!<�M7�U�H�a��!���|��,QI��?�%����k�Cy�]�����$�O��qĸiLhPS���$?��eҲQh�{%꒜�W�q8�(%��]���}���jG�c7HvV�+u��_P?���-�l�|�1�a��l��epfvnh6�rY����潏�J�g`�Gx�k���֚����a[�k��Ǘ^��r�N���z8'�G����1������મ���t�K�e2Η��T3��@�e0��
�J����	���Q,סn��r�vi�ӥ��'(��k��<8��]�E��W���:W�)Œ�qZ�ה������${C_De�쮜�"{6�U���u�����,�A�?B:$Ĕ�p��h�K��,K����:�>�H=izǀi��HWԜ@���`��=��/�v�8��
õ�g�*I�e���S��dx��}�����訒Q�AN;3҄(��_��-���W�t�F�m��p���$À�Gf�F�:X��-L����u�zP�?�S�Ԥ5���o� �2"�"5L�#���́cȆzC��w�Q������G~�����%�_n��
"W�o�-;���@~��G0c���hkc#ۃ�n#���E��O�q�R�v$ޮ���}WK��f�L����ӬJC���B	0eMd����H?�m~��-r<@l��sf�Bn���tE���Z�evu!Ԩ������_�*�b-�jf�����ȄQ���P���>����.BA\�>����9��w?��%��E[�v_VOE1<����8[��Μ�f�D���^���l?'ލ~�v��OS�k�n��9C�A����ϳ�n�֘Q�m �:k�y����A�N/�^�k�$>!`Q��q�!���w��h�ZJ����CO��q�O��[���r�c|Y*]]d�+�(�N���ȉ��2�PPMN������J�[�#&<���InXE7m+�HQ���ʈӥз	V�G<��ӽhU�E�����o�˝�9'�+ם��!���1��n�RV�L�.�Y��q��9u��&-���s�AW9T�S�����'	\A��x��*��y���q��V)8���e)v��v�M��_I���-�i&�_)|N�4���L�˶,.Vq�2��|�ѐu��fX9^�.;�aIT!�w�ܛ�J�ׯ��I�u�_��N&�_/+���pX-w������Pp��vb�d�q���
��O%e��Ɋ�����ҭW�� 1���C=-���	��Jd�"C�Ď߅9t;	���U{��=�A�1�L�޲T\��X
/M���s�۝�ix��D�T����l1��RV|�f�nZ����T�S�t3yp��|ݩ(V��]���ʮTj`�~G���/A�?e&mt��r��H��B���`�!S��*J�x�:鱋7�=�=_�vK'Ӑ�6�i���ЖZٰGa��L]���҉0��1��H*XW�����������ك��e��e��O�qLJ4t 䱕$V��O���k���=�l��R����#�� �����ײ?�գ	�;~��	L�7��$�\�K�Z	Ň����Y���TZ���<��<jN��*���a_uAL���4qچɒ��ύ�)���:�FT����� �+�^gʯP�a3�m��w$J�s��#a z0+���bB����48�I�]����M����cG6�b{, ��t�FO� _W瓝�����A�HGcMS�銻=G��|�-�#H��3s�znkS��'�<?�j{��^�t���ͣ&���޸m�a��'4�y�]5�(��A�yf��T1�9U85k�=��C�B�ÙmF�<�"����U����Sa����N���d����e6Kpkb�|i��?�sB	�bi�A���;�'��稂ƒc�t������K�TYf��T��%��ƣ�x�x��P�	7� �g����F8!�ٖ|�8���sgLq�9�/�?���1��R#lW���rFq����眵��&&-��U�������h#�85S[�*�Q�Y�c�!�%ei�����:5{aƳ��^�v�P�f�:xü�Gwt�Z�
�̾B��`��(�����u�M�NYӃ���^CM-� �`nn8��Q�U�H_��~�p)&/�q?M�eR�YY�WX��O%ج=�U�����m��,���76��射ȪG��%H���T͌M�0���J���o=����(P�yj�y���~�D�pz�f�.��6J ̠�  @�,.�ڸ�G#�~k��1�h���'3�yG���ͽ��xo%��ar.�?ޢ��~���t5�s����[�,�����ѩ�~����#ҽ�>�<pz`��9�o���u�T b� QQ�Jxvi�E[��@�������6�*�xr5,u���u�&��LD�	3n�� ��Y�?�sq����"n�3�a6���F/[<��DI(��6�����sm���+��¥Z�������ᆶ����)����W�9���,�96�1Sݾ�1���'o��&Y�k��p\�{��p<n@"qC��¼��7���H��[՜�ׂ�����cN�?L��k�q��OQ�)���$y�g�.��!i��w���ˋZ��/�,z�&�/Y�Y��_�c�;��`;��5<�A��RہH'yV���W"�΀0�A��rކ6�3����}+�c��hW��	�/�;1O �6P�80���C^�����z�"gMz�b�1��]�C4&���o�$/�y�	[@hx�'��9hZS��>P���L��-�ʯ�}�������~����M��������)�Gtq@w�q�	� �xs=�M/Ƶ�_|��]�+\va̖7����j�3�����)�����kq��1������BG>v�e;3��㽿�����V�y�2|�����bw��P��~���Ez��[= �]��W�p���=���=�H��J������i�ú���{��K^�ק@�9�$�7���pl^0����5y��T��^e�o4p��0t.��ģIV��L���E�*�'�#�T��ǧ��ķ�zX�o�I��WG�W�G�b+s�'�U���M]u��@�kx�Ep�@oMK���ML᎜��N�̼�))>��v���%���L%2�����8;�A��$��q�O[Fo�\%�Q�F���w��.7�
/
�#�IvWQ�pO�� w�lAp�\�.�f����QD���<�h��a�`��C3C��1o�4�z��nh8J�
&6# �z�}|��P �����0`��?�{1�i�vkË���]�b�*;|:Ɯ��ќ;�Ԏ��	e	�����1fu�?�)�5 U�V�/�QX����f�YhW�fڇ�*����ۧ�v
.D}e�ҾI)u0�g�I�S��U"���v�����B��	
�@�v%���}�E%�0���j�N��Qх�%�����ݴ�����Gq����YA�X��ؒ�]H��5���,�Z<������;��,s�����U�����]����ꡦ��L8�*l�,����#n�������ٷ��6�BB]�Wb|���Z�Y��p�p䠏�j��A�T�_5��ܱ�̣s��[�}�Fx���*�-�NZ�k���d�Ġִ_/L�����P��Ҥ�����T��B��b�����e؃��E��K=�2E��I��sK��6
��>�Y�ѣ̕Js���yV_M�k;���0�M�Q��;'R;}뮲�2um�)d~�$G{��������v�`"T�d�mđ�;܁1��M�p��]���`�!�jH����r���Z2W>�;x����3ƥ�TJ���9n>��G0�S�%��8c��5���u����s2����C�]��-⟈�e�ͦ�àhJڨ���^����kh��{�n�|��0�%��iL{�	r�f�`���heWa�N�$�ػh�	�i-@�m��)R��}'��ZZx���=�{G�v�v�N�X����J����F�	���F��E�����V���#"���c�c��
OB97���tF�����%f�8��L4]X�^��7�7
q�;w#�-xwu��n�}�U<��+��"�1�E%y&��Qӂ�Z���^���`��Z2��ψx��Xl:_����B��I��f��}�pT�M��h<�+	Hx�0e�Z������S{c?�{W��i���ˁ�
:�{�����25]�Ը3ʲ ��7ֳI�E����~��س�u9�d/�5����qE����γA�'��h�Cd#p�E��N���N���װaG��V�!�,��G*t���_L��j���t(M.�KW�N�M���]RPp�P�D����z\%G�|���G��k&8�][�{��K0�h2�8!n:qAre�0������/����I-�E���}������9�@7^�a��l8�FY�/GϜt�,�g�@0ٛ��|q6Zӷv�K=�P"��%��;x����QBRw�>i��A#��O�'�+����T"%`n�&L6m�9)7���b�sE�b&<��:?jx=*�|q`x��4��<���-��Ovp�K�h3��Ӫ�s|��
:�Vp|�x���U�Bd�;�݁c��X��u_">�1vg��"MqV�z�!�{dHQ�K�yEĶ��Hx�$�nkQ�qO�X��g�4إB4�%Ʀ�rO�M�鋃|�k���u8ޥ� ���	+h���7kS#�Lԅ�$��Rl�Qw�_|��:�T��pǺ����h=p��0?=9���<�Áކ��V�\�?o��~���&V��^P#�ܘ��@��e)sb6���p�${����6��B��)��x�������zo��.����	>7�)�ۮU�qiŕ#:f�C,�C�[��h����eo 8�S�۪��{�����̕����Iv��ܫZ�Ns4K{V��\�lm�Q{�>���2�����o�N����?u��X��ИC�W���e>������ſ���ϕ������!GP.q@.>�v�Ͷ��:�Y"�	���j�3k,��n��UF�Iu��x�`ѹ���>K�P
��8�&���h�h'S(���(�qsKJ�-B�K�7:���0��j'�����8��ul�;X�^u�hM�r��l|��E��!�	*� �h�X�v��1���H��*��4���P<j�i�=�t�Z~j �@f6\�<sW�H��j��׼oj���1�N<�j�7��`���7�W��)��G�u{�l��ٷK�<}��#��eZvˎ�12�]k�{�C��O�;�.��K��hՙ�0��E~gO��x����2��!S@�L�@�j.(,^�$t������݉����p�\Z���#��7rV�Y- �|�h���L(?AC�WO"������*�ݿ���Y�9���B�����j�D���d$	�
�'YT:2Eq�f.'���
T�M�f����J�2�Wld���X׬yYKP	0^^Ε��宿\S˱���߃��O�^I	�=�}h&Z�aU3k�W��Ȇ,v-sM�v�`�+|�]� �R_d��� �*�"g��� I��Fw��By���~�B��ɪ��?��N��G3�_�&�������ߍB�֢�O��oI�ܟ>��&�z~D^&����!@��`-��E�� �u�O�]������4�-f�;&���]�^�_qe3
o2�˴�̋I��z�յz;Qi�lA���Q���%PW�=81%*8cp�E��UaL����rW��'?�aoT77��Â}�$>���@i��Hj�&�+���@Q�z-�_��g}���e�ntm��R�W����;DU�� �L�Ew7�/I�LC������K�@�yţ��u���W������y��&s|e �z�Sz^��`��{��,�u������CBc�W���/cE�cb�RNf��D��%�{. 1���PG"���oʌ��z��J�䄋��N^ú�7��G��
<u3�����2b���	�kh(�CqX���Vi۩��Y�>��n�!	`��̡���`��S�i�����r �u�z�8��}}��s�968U�R����[֫n�K��G��O4�Hܕ�Ft�ٟ�Ȗ�w(�Ч��YOL�mb��(�4y�[�P���ݚ+�3�ט��fΝ�n�w��sT�d<6$��I?o�R��S�C7{�� �=![���}��R\QE��K1.ԳM�7�=v�e��e�s�N�o�e��%�Z����>�Ȥjݼ��i|%'=*�M�'�=�N�ȴubp��/7@�>�0 qI�V��t�z1d#��$,y(N@ҊK؟;F%���<=�}Q�nz��|����[���*�ċ���9D�R	�0{ ��� gDXWu�.�c��h�{H#ᴺ[A�`�-��r�	���xF=�]��9�h�	X-�i�p�y��(��<�=�cOrD��a�%")x�V�ǎjYp������W�n�2�r��t�"A�p�����/�`�o(���2�N	� ���zX�����QM��V�\=��_oL��w�p�ޗ�C�7��	B�@�����p>h��@�h���J �f�1l9p7QWS�nH���ڿ�4�d��h����Ir"!��ʿ�&L�Ϡ@�>��1a����htx�"!;|-7)��:��54���uP⫻��v=��8�b@	���K����n>�̥�VP�4'
��e��~W6H��;�L����%���8��n�������;��b(�n��DPS��撃"�_�<iU�Q2�¼�d�tG�Ig��[�=�1G�� ���"
h:�<ӭ��"�C�z��1��0 w]&-�8A���1����=�h �[f���"r���񿼭!���O���?T,8�%t�e��3�tJ?�B�??ngj�M(��ˀEp�Ғ���>Er�(�Vc��<�]�&�X�ZE�� gz3�~c?lg�歃�f��k�l���nb�3{ R�����,�VB?�饺����������z'�U.~{�H �Y��*FE|:��M6��*�	g����h�_"�H�æߟרݏ+gЃM�(8!l3謑��+�ϴcH�S��q)�>�������-i�Ѱ������o��
�!�#�[4�k��l��>vk0�JF:m�'{�Z�fH������6s��5�{慄�m�񝠹��nfl�;+c�u��7W��c{	��͇d�e2�8��s�7��S@z���Eʹ�;�u&��UD}�a����M�8jwR�`�]�X�C>�V��X�0��%�M��=���搅���Ll�����y�(W�*�3���v'ǩ���x9��/�c*�Y��B|��<e��/�(��P��,C��A]�4Z�%��1�|>A�{�U�W���֧��H�����b-�	��Ky�Jb�hꙈ��F�v�ҝ䧯N�Y��ޞ�D��\h�Ns�����Ľ}/�w,BW�P���ap�qi�Ǆ{�gY�~�� ��	�%�Мר����`�Rܬz�Q�B�y�X&�w�К�"��V�~��5aN�N���� ��9�_"E��|���;k��R�G*;>��:N�����
{+�����`it)6~-.K��l��Ք��t�iۡ���zt}�'�X3��C��B��׮˛�ĤYٶ��S�Q� fD���8@h�������?��>T���nx��o^o9t����M�����K���̝&R	�V=�ΓLGh��Lwv��A*��oVA�=��0�n,R����Q��[��χ{Ϸ%L�!?<���θ��߆a�F/�^��i</")�F�-M[�%r	IM\�E�h+kC<P��u�<V�3n������I�^ós��X�#8�%��&
;	�t��%���Z�j���-��~a`Z�*�ɖ^l�&�������'=�(č%���F���%|�nꊹ�/RtL�#*T:��y����̦:A�Xjџ�����`uw������.թ�hl��T�B�������Ʉ���z�;��'�o�Md)*����o���7c_�Qϰ�<�klid��4N�X�~�C��i0��1Ff穿�4p�Ԋ=�|�jV�D����O�����-���Y#�QC�R�����j,��~�%|\YF5�N�Yԍz3%^�br ���&Op��t��^9�s}8PǛ���2�^>��h�ڱ����s�ۗ�\2"̸ۙ�����2B�ŗ�p����.��D�ό4�3 ��zY�'3HŨI8�-�K*-࿲�O{2m��ߞ�	�C�	��Hx�EV(āqg-�a�⨉�η�^���u^_��"���+[K�^ʋ�z%�)��L}+~�Q��ҫ�[L����]|:�H���Vr� ff�1�9�H��d
P`[���[S9k�?�h���s|)s��JM޲�<���gpV�T��
+��V��M{�)&�1r�$�����j��OB��.��۸/�����Ҫ6� y��[��=�P,#���,�p�*�k��ifY�����SW��c���fM��� � �7e�ȍ�L�dq�4D,�j�����v��uJ�faQy��.ѕ'�(�ן��a��҇�(i2������t�k�lYg�i�aV��㘥"��S:F���OR�)F���`�{�W�eȰyq��jZ������z�7��#1pj8��o��Wy=;���K$��-��07�H���*����s�I���_���� ���Ōo$�0�T��ِP�ܸ 0��-��T�rͪB��^5����"r�]��UN�/x���L�Ah�٩�t��XvE9�*m_up2��k�0���C(S�Q&��aֽ煨S �pw>�|Ѵ��hcd~�#�,I`DG�2��[&�"yFp���i����ߐ*��l����[�������o���}Ej��f��i��AB��)wu��V��;�����J2�
��ZA����{*B܍�M�X2��E�5'Đc��+7�;:fW��R@U�=��&@�7����-s�}ƌ�UG�=�8c���о
�C$=jf�D-d8�[�Q$��;ϥ���[6�~L�h# ��+����VѨS�Fa��M�qߊ�Ez��i����5�DG��,~!�
p�ڛ�������$|VK�a�X����kϓ�3`3t�y�̯��\$��f�g��I�V��=�=���������f����h@�q\�mD�{�L���@M�2�ƌ�h��$WE�\�V7��'X@��L[���|ؠ��[}#�`�)�߿�i���:^z7�ޛ�~$��$U�p��kdv�q���La����$[_(�9�f�NY)ٯr5�+��K:�2jm�^N��z-S�f٧���*p{=l�@���\Mi������N��!�� M�v_&�p,�#[C���&�jʰ����D߾���Ov v���"}�5��U��1W�m�;֕\K��g C�=�6�GC�- ��h�Q)-\����M�-&?�3��2�3+s�@k�D�;��e?�U�Q�e�+y�(&С�%^�1��EhoG����{��I]��Z����l:���18RI|�����J��R��4�W��䆽�x�Zٽr�Û���}�b�I[�#%��L2�C�*��䶀�hs�a~�?\�����B6�7ڋ�X� yT��@� �1�[��3�}:�@��SAyF<�^���~��>Z
`vEAr�Nf:�q�V�H��Ƿ��쥁��`g���V~�R����̙�
��L<fRE��Mz����5��P� �٪�H���o�:^��4߳�x������F�3�
��/��[�K����N��N������I��j2:c�X5���~�#,�q�c�Q�Nɍfw:ggkM'	�m��u��yK�IS1��*����{o�.:V�r��q�
@�zl�� �`OVh]���V�,��{����7��.��6��@� �`��FKV~��]��:���B��dOk�R.�뚂���B��X|d�0a�x�C���{��y�hE�F������ �'�-��w�ͫ�����)` <�}�1��J�Nr��Q�\M����g��B��R͋MCs<���Ռ�C��D#����p�sc��f�c�O�!t��\.K�\��00�W(m|q�5�D�Q��c�{i�Z9��#�a	��m}�a[V�8uDC,I����܇�|E,j���ƙ?0�B~�(\]���^��::�1�=�-f��[
@�,]�^�b�P����ѭ^�?/�]K3GA�Z��ё�o�������6oƟ�����#���G07pC�UX��
�`��S(�&r�'g�����jI�hY����5f�۶kZi��|�FA��ȶC��_��<�e�K��V����Ԋ�F�;�hO sk�uiK��ܢn�c9��3��� ��0)�K��z��8H����Hu��~��Ɛ����e� �N.i��%{����X��aGW)��(�r����y��8�<ߏ��?>�5W��	Z�o������B˒:��'�+����[�/���I�g�'��`�9�=��Z��bE���qվ���s#%�����\���[���Xt�}�Kf�:~�~�!}g���ۚ����χ@OZ?�cF��i��̊���r5�mOwx��	��h�[�5�E8�d�f�圏����9a!�r�M3�]m�����%%hm^y����K�]���a3�����⢻u�->�sa`?D�/C����4�^,s���.�}���a�<��ښJ�?a��e�t]G+˒�=����&ѡ��"On"ɫUe= �H�LL*���Y]W`G�W�򋼒�ұX���b2��!���')X���N8�%�(:л�Eeu�`��#���T)��LA�b���y�t��̮΁�	�����Ar��̨G�\�M>��o4^:����I T�6�i)0)M��M����Sqm�^�К�/�_��L+a3��$��q-oJw���ƴ�A7����e��H�Wqa4��ao�E+�D7�2�ֻXgd����Z��R�9�4��J'������x!|-^�'$�(�Z�=G