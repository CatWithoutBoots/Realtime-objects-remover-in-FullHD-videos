��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�Pk���<�T2���݉�a��<�B�t�7$@�}��K#L!9p��ud��^ڵ�@j��Ff{�緄��@~�z���G*FIC�����J�S0��
j�xp�M�,���*_��:h8Y��E���V-�y���(�wG�:G;����l{h-�9&�Q�/1��Dz�3�� 	�.�؅D1��4��7;��50�S�'�i7�Ҕ!Ԭ��A��L���܆?���j0y7GD�o�֫/-�\����D�u�X@���s�5�#nN���2��ǂ�u� �l"S")���� �J�8OI�# ����t����C$mzi<�efph��sA��O�C��
:�> �WTS���S�GZ��>-6����-⪹ZR��<��~��I<N0X�2c�2��|5�$Y�in�q�>���bR+�%�
���)�e؃ $rw��|��c���];;NB�/Wϲ��Րq�A��?��SCN�Lt�.�n���rQ��0����|��٨���0�����/T�6�+�bgO�t�<b����J9���Lq�
R��	;�>8�_`n�hF|l�
e��#��˜�_�B�(��k����ǀl��W�Պ@�?BTZ��w��[Dg�M��r?�qj4�����6"�G�<�T�W�҂C���U7�oi6NZ����e�x'7�$ۯ�'9�P�_&ʴޢk/'��[~i��P�v��_A{8,�ǄKa�ԁ p���nq�T�B7$��U�U~C���W ��p�E��q��]E2{	�>��~��~$�%1���d 䢱�Dw`POg����C�1NW�t tڻ������� ����_�'.��o?��qBq�D�o&��F/c6�=�z�M�p�݊��u�}G�	Rvse[ �����(�����-cƿZ;`u�/`A��cb�G)i�Z�6=G�]�&S�B�(7�I�c��o��S&>�7̃Қ�E�����Ok&駆�ti�zol�V_��=�҈��C�8-t��9i���Z�&X�\�/�λ��1��
r�n���J�+��f�S�TXDv���G<�o��)ո������<��A��'L��PAt�z��2����W(�~����n��\��Ƌ �3TZL@�<�Kg��ykXZ��aBL�R��j�}7Ha�,r�5����P1�I�nR����bP9�.�K$�)0Z����w)��z�K�/�+�`븸�����R��*�ej��!0�<IC��)�E��4�'�Ș���B���66P��^	E�䜶���g�v�l{�2����c�)-�!�s��}d�:5,_�ew<��u�Ŝc;.ZG@�T�m�(%�Jy{��+d�<����@���U3�>���$H�������j����%��y\������σ8&Vy2����\U(�����>��P���{������06p���P��H�����lSaf��#�S���(]�Hʃg�0�B���~�\�;m� D�uh���bns��s���qC�kaR�g=���P�q��<����WD�+k�PF�-��9`��N��+�[ÒY_�	����Dt���.��>���@��򅁊k�>Q����m�C 4]��P����'I�t�8��+�8le�]`U�qS�i:�b�t������X�.\�ã(�n �����"�p�kٌ���.�T�T��2�z��q�D�!ʐ�2TT�b>�Jʄ�?ӓ��]+�Y6�K�j蝏o�����#joQ�68nH{˕Qa��C���W������|��$��u@���¹��\:��W��G����֨��B-3�ܔP�u�C�&J�V��th@){�#?��5����{�4kSTr~<�\���2���S{T�a�R�m f�� ���<���:�R �(�`)���c"�ކ��<`����b�6�Q5���*�MSzMf���~ �6#�>&*ȱ䧾8�T����9&�u��y$���Z�0� ��Xj������͔2���H�*���>eL_��5�D�_.�d�#��f'I�6��I�/\��#$��ؽ��>A<��Lw�"	�L�-�}A�V_���({>�.��Be�5/��:<�?	�� �o��xDĚY];9@Y�L�av��H�3(�nM0_5�@a��&�4MFp�٧�Źj��8�"�,if	�����x!�_^in��w {4��n�9F?n'&FGJ�!��gA��LV��~�9Hp��f'�'�?{0j��W]i�p�wݬ� 8��~�Z��@/�vO�{�p���J������XKp\���t�) �����֝&�Uq��o�9��f��˩�����MUӷ����@	��+`��pPݭYK����;��T��������jG��k��J����}��D[�cB��6>/�i��i���|��R2$���̎;�XmHM<'�fՎ�=t��|$k���M���ԗ,�J&&魧4G1���yev�}�S����F���
�D�8ǖ򃏃⣓)��31y^Q�q��a#c���C���؊���j+"gO��/��Yi�*��)z+�G�'�ޤ����5�{{J^�r�qԫԲ��S�|t|,����S�t�4{�Ӊ�$�|�n���%��h���c��_����)k և6dn�r��{5�2��'`ALx%�(���-�}�����ؑ���:� �L����&��� ZQ����,��:�����A�%3k� ����	թ=��Xc9<ʷ���㎖ɸx�����7�� �"��:R=�Q�<�����>N��Bp1҄|ꪗ�o��{�?�0�^l���ۀe�^`�i�c��sU��*q��Zb}��1�&�ށ+Fc�8�[�v>��+�e¨�V�syR)������ߓ�����5�:e���=Y��(3o��Ϩ!�z��bȭ�a��c1YY���z��G��m�*����+.���cq!z�>�1��W
ۆ���.b9�g�_H�^�Y��Z�}Y.��b��Hn�ʎ��z*��7v���j���������쵝�}���W6]���d�t��A =,�3�����onN�V�w�Pir���r�Gd��>W�c֯.������p�� cl��~�h{G�`�Â�['C�CM�<�3mL�,��,��i�p)�R���C�|+j�&.E�,�r/���D`�oF9�)�+��W���fD��}T�×�1����	�)`Hࠢ����g�LY�@I(���D���[�q��5~�K��4 ��������O+M�����8"�;��x3����W>��u��_����� yA[Ƅ@�_@�9��E{��}�ɭ�|�+R���Qɇ2i���.��%��z��􍭬<ױ�tX<$�����BB�G�,	��.v�C����~��&h��
���me�q����XC�=���j���8�s)
p5���sv E�NR��۲����Y���T���f�6U�>��Uu��6b�h���ػ�&G�����,ˏ��yVѕ���������_�+�3��G����];૽��tòg̋�I���P��ϩ�t< ��������M+��/�j�i��ob�����宔'Wb�bCDP��!��'�*<hp@G8�J:+u=��g���,���G_9��+�Otvoq���A�@B�ĲZ!�O��;r��f�&๬�����TD��vD��8W۫r��J��&���$]�ɇ~����pg�j=�D�"x�DK@��J�����1g��6THy'���q�-�GP-�^��b3�.��C8�@�������@�.���dO婀�f��d4>O�Ƹ�6�a�U<���^��D}fN۵��_��Ƥw���@�!�<Y���:~�y�OH�3D�X;:���Ri���u+��ن��u��	�ג����7��e�#J��L�,�fL|D#�~�_�����Ah���ID�HD����� OE�� È�˭�X��MO�_x�@XxyQ^P�ÂcX�~�N�`��ೇ1y��+��[O�L�>���q�8׸��c�b~�)��>ґ{��X��nO~p�K�L���Y)m�����w�c8DK.�	�&���������+vv.&��b9�@�Ƿ��������:=��(�׶И����Z�	f�؄ٲ&�_X��]Lm����:����C�6�������K�!�j�13����9/)o�6x����t��;��a�ЕxR�s)�+��b�w�p�'�x_�d�j��Q:�?��<H�Y�(�v>~)���&��w!,�0�<n4gPmľa��Y�M��@o*����w][��T�!�Wl5�����w�Ld��6a9u+ޣ�2xt�k�}j����`�,��Wm�y֨�%�a��h��0t<IѺW�Z�:�J�Fu���>Dw4#zA�;t����%L�����@�V��z���|û)e�:&���l�&-x����~���T@�L��;pS=i���+��#����������r$���O��@���_�*���8�S���!R��j]��y�>Ń�>.��\�1��H"�0�M��W ��haU0����[���23��������N���AW�17��:x9>����>���Oܻ/�0a��V�w���%�y\������{�<ȱ���C%�����i�<;ƚMkԙ`�0��=)_^\�-3�v�!1��l��5�CE:s��N��5��2��v�P2�*`�R�����X߿60 .��<-��������mj	9_-3�ɽ3�^�!�d��9rjS��Ң��KGj�?ק"Pnr�=:�]�׈����Vd���>�m�.M�7玸46&��$O9�s�1Y0������enm�f���M�r�:>�;@���M������'�MZ�ܺ�v@C�(�@]w
e�}���D��P^A6���oء�z��C$��
���I���G~D#�f���L���;�E�|��nv�&�FO{T!�~��y�d&l��%;�_ +����Yޭ��e4��N�e�1݈�r�(0���@��}���*.KS�H��O�4ɉ��nS_"�[(Sp.�����"�2S�<z�W�q��_5i%�d�{�eTcQ��*>V�`]��,T*j�
�N����Tj�[<�K��MS��s�ͦ��R��:.~�����Z��2Y	�F ��{��f"Fd���-M�g��Th��y:��J2#�Gt�ڼ����[��Д�H܇�#ʏ�-7�}���.w��9@?�r4�ؑ��l]V�� �OWJXTF#��y�Ώ8�
���9�����)����Ho��\�����7��
]a�6��3y�%�9"�@J`7��� ����v����^�(۩=/���!MA%�A��a���<��?`tƓ���s/��aIԊ|[�,��@��N�8}�o����:ꇦ��]��A�>�K0�H�<�,��px��S}K}m�sv�
�ީ��Z˙��M������p�z>n,;�x���E�B�Ib-eG�0����⋱���i�s^7�@�f8(���{�_b$�8'�����#ح�����X ���g7)�^Ú#�����}V\뎮�Vu��Zy��1G�#+��ŭ�;7!=��^h�a�@�[i�v�n��܃�q����0��y���q��Q����Y�7*�j���l/���#��a��{�	��c1�?Ë��吓���2A�) �a�y���8�Rk��,��PYe}F8�T�˾Þ+,,>�ra�L=�<��	N����
C�����5E'a"IOsH"����� c��	o��Z�`b�]�@��j'�4*@�ǐ�R1���_�W�q�s,rjHT�'���g©�?�ٻ�������W.MTn_YZj?�5��Ŀ�V	�rǒ����Q�l�(���T�k��'��Z?��=�b�a���.���G�^�<��7����N�f�V2s�;�-��2�gDے��QPMŦ���b��+?(!�6.yF�����0�h 
`x1�[��K'(�$Q�W[���s��|����n�u�kwP�Cm�4ӥ��-���tk[8Is0)+-�v p�[�;�����q�UU���uj��¥�1�Z{ì��H�%���T�*�g?�륨%Fb����x
=������6?2��3�������ڳ)T���(ڣ�6rw�H�_{d��
t���h<���
�b�,z!�R��"��Ǐ��J�(v+2H�B����'H�k\��8�����aL��fVx��$C#�������^Y�D�x�������[SתJ׶" �*�B4�=)�����t�.R㕠nRW���H�q�X���39[���J�lq����.���󈴫�Q��z���/47�����&��m��; �OxM|��Ϻ�Xak��j�3��d�G��nt�'8A���P6�\c�b�C1~�:��X�������CAN��/e!4��珅��9V�1����ʚ:�!��`��|C$��S���e"|�C{�=z�>h��	��X�n�m������{>�R����dyD�������0���%��}e=���M��9΍Y0��\K�SV�Y4��h�LdV��e�:���'J���88���'��+�j��<x��q���G Q�� ��q �˱β~�a�k�O8X�U��n�%ɠ����^�Q�s�z��J�tƤ�
��(R��9~:�N��<�"�ZtD��#���8���N�p'v�������;1\,Cΐ�T����Ya娧,��~-��o���� �:����������*�`�ې��������� �'3�҅>{mGJ?Hv��E-<�Y�O��7M{H�;�^��Dl�/������Wu��x=�fO�2Mq!W�4�^����"����\}7-�Y�_���@$���#���e�i/���-�om�m�c_\X��蚇�+�N�v�m��vG"cPU�>�ol���ߝ��,�r�?=����x��+2�"Ւ-�A{ �x�5���}��=r�s�WS�Pխ��u�ݐp����'q��Y�"�a����GӁ���=g*ś�M�V�����"�6��D<j-���z��7�07��z�k�J�{f,UDF�C��H�o�C7/��Z�Zk���_�P��	�E�}h���Z��L����4���^]!�����;)�j�ȧ=��k)�V����N6����~"��5�?��!���5OWt��l-)Fe �~tu�I�i9��5����'����I���r	^p�[�1ď���ޤ��ZS�)����r�L���qUN�cr�D�"������>��~���4u��մ/e��V������96�y�eUa�G=ﱂ[����q�zo���s7�w'�����Aj��|����>�ĕV��>:I��z�M��Tg��74Yeܙ��� C�d��2�:ߍ~�!�ޥ�5g��~�p��p4��+���Z/G�����cq:)*�arq����Nڢ��=X���@�V�~AW�g(�$��>���[o�l��HGڄ>��xz*�X�X�i�E_�����3�E��^�3Gϙ��$^f��Ѱ�]�+j3�_� �]`T��嘐{�)��;/*97m��S���Y�_���}B���P��i��N� �P�ۆ�}G8�T���0��;�ŸsM�CK�B��I�gr��_7틎����W<i�K����y��3Jq_틝��OX�1A8٬k�l�jR�hl��G�����j�^��b��3���K�q�_��#����v" �.U���T�n�|�d���A&�L�^z0�yA�$|\�߂����+�1�ȍ�1�=�y� Jظ礰{��GN�M�������G�2����C�(#�� ��j����a�Q�~_���� ��i�c�K�|Tu�*������JG3:|�U�ۉQ���v�y��%9V�p3@?Җ�9"pځ
��0Mjyg�~�	�r>o�~�q��C�73Ӱ��Ķ��ep���(���/;���/;�(�:`b�������-o�+�2	z�MhG�a=��VSc�Fȿ���nd��N;�@N�_��LؿWd�CQO9-_>Yu8W��z:l�%��⌢�� ���{�D$w�v��'�Fm�oJd*j������f�`wb����7I�����"�I�flD{R���%��sX��̞�3Q��^k����X�]~�R�rKc���?o��;|�>�X��J:��]߹�ڲ\}?�r��}�����ܲ.|���Y�)_��O�M��[��k�l�T{J���8f�Se����&HO�+��ҨwMz��ŠD�ī�I�C�z��9�Cږ��ЊM���[꤀�I���)p�.�Aq�jH%�{�D��k��u��3h)PS]�x:��B��sԣo�� ��>�4(i�p�j��AQ�}�m�q�>a��R�u-���V:����-P̠F�/�|fޗ�8R�WV��b;c3@���X�
�eͿ�Z�=L�4��K�����.
'��6a"o����I����ÂG�|�C��&)Y�F�_��"�)�ؓ�T���c����7��YE��;�ц!ѧt.q_�]H)�]����oR���홱�ݛ:�l�Rō���&�7�b���e�q��¥Q���U�����R��S'���r���g��>�+����l-=+��c���shA<�"�-1J(��ɶG�G��^�c����|�2���f�� 5FK,�#�|?�]�m;?�����%&{��,F��������fh��f)*'�cɚm̀F�6�+���z�ᢲA�>J����IN��}��W{42W&zAk����+"��mC/<�NP@�H��HD&��a�^pQ[�Ͷ|�e3J�}��_��b��:A/ ���f.��ȼt���ذX�ov�rV�ƞzE�H�_��R���O�x�0�n�kDn�E;��I��gS�6=��q�-��l+VQ�/��읨�u�*�7j��Z'%�zd�J�A��M�T��� ��CL��l��%_��&��s�~����%�j�]{���)�n��[��M<��_٥|�)K �V&�4<F��%�n��q�E��Vr��h��P�`�\-K�
/��ʄz]���yj�ܞ���o��j���^��n%��;��v?m�wF����"8NC�`��,��qI�{ܺ�P����Z{�18�F�,*�xtLbV��='E����5���~��`�>1�]�VP#�u�q���E�ӵ�Z����؏x�<���*���'�;t�+�ު�4�\O��δ먈s�����\�A,/Sf��:�T�����i%��#g���#�J�)�!�����u��������DUB�Hu1��K#�3�	�����2�$��Wi乾��W7���[R�����)ؽ~����u�a�
x��B�@�21  ];%i˩�������%��G���G�i��i��,�b�hF{8���!&�`n���i߸L�y�Y�R5YC2V����xM08��,��0�P5/ӹ|
y`SEq�KD1�6���n�5��X�t&� X$DI�RQ�s|v��u1 �[���+�;ګ/��X|�yΫu-�� �;-��2�{X�����U\hD����}����
n$�!�Ox�w���L��Z��� R�����]�T�TfJ��Hr&�+�"c�X8��n��/��#�%�A��/�hOy���Rqğ;�B�>�Z(Ѥ����wL�s��HK���3cj���^u�9`�f+n��,H�9�B_�"�L��~��&z�!(�=W2�6�!�^7��.!�1O�5A�Ζ.�597�Us���bXR�c,�1����s��6��R�k���$������ւ	\Sn����޼ʠ�|Y�{�6����I��9��U�Y�&P���{�c&U���[���M��UqL��x!�p�cp��(x��Eح0�Ye����!9#��S���_ST���\::���Cx'�&���|)��ɃB�nI�"::��ҵ���hz�X�<8������q��A"�伻@��x�G,6'��^������I!;��{T��ď�p��N�#�{5�4�n�e#��Y��#l�{Q�¾3��u7H\�}xSx�%���
���U��4���]�_��യB�ϻ���nH����d�z�5�XG�${�43\dqǢ� ��K��(����M��ME�Ȼu����Ǟ�Ƅ*����E�zu#�����t�8
ow�yNt�4ln��Dc�������I{�ʞR�i߼��8��V���.s]��Ι�kG��x��t���3��ƅnc�Z��(�E�E�ti;�����n͊�L��5��$����B)���|~2ο����4���婗M�g���nF ����(�o�$8�p\ [��SqǦݬZ�o��S-i��ۑTg�qş�,�8˞Z�j���:��s��X!RI')�9S�"���O�ݸ�C�<Z�̃�){�ޕ$ZK*+���u��uhpM��x���B��\:b��Juy#��4th�ʈw�Ӫ�*	����Ɩ<���NΪ0b��n���I���6��ڽbH'�4:U����ǚ��أp7_n��!�5}?�[��K�x�`�VW��'Ȕ\"�����Cߪ�' �Y�Zڭ�Xn@��\O��.�%��UڜFE��HܘyZ�0�vF蜹�h�A*g�e�&��ǇfD�*/�F����J�Te��%~��h3aZ�s�(��3��w��VE[��x/T���F�2bEr�C
���O�5�8~��Yv ��G���f�1U윮$`�P/:2�rM��2��h�w���;I3-�s�P�@9P����&/�'}NӘJt=�I�/�NS��-%���֖5��店C)���7��M�'юu������S��VH$����4�4H�h�iu�j���D]B��K%������(�0[̤�~7�mZ.]��a/a����R�i����\�wXL�0i���(/�ZA�2�6Jr3�P�:��pf��J�il'tc���9��P5?R��C��R瘇��l�dIr(��!�s8���^!�_�6�\9UH쵕m��AJWK\���;[VM����v�	;���"�ɂ%��5��Ŀ�g.��P��"�u�Q��,~��}�J�Dk�ۄ䯛�tG��h.rҖIE5�o���W�8y���|dx��J��H?!��ك����!`��a�r^\�k`��h$x�^fL?^߆\�~���ww�a���V��UUf��6aL摾�%%��J�7���Ϙs@��*�w}���[��-ԥK���]�v��S��]7lA]"�����������W�a�L�a���
�n6G�3Jo���;J��Q��9�nC�KGI�s����x��j�Bhf˭}X,<s��т+ɡk�2قW((��/�=-�F�B���3�f�#ItBTM��dX��
0��������ձ���If����fj���E��Ӯ�eX�BpT�"J�"Ю��@�h���@��n_�h��q!	66Ut$ηCB�ܐ�Hmf����C�Co7�a����/YzC�?*���L�+�c^�q�R���Ж��-���X6�<%����2i��0��uU�z�����h� �`��ׁ>౶�xq�D���Ǳ���i��i܊���bnzcud_ꢮ׏v��:����gpv���v�ִ��g��c$ܪ���e7��Y�_R�uG��J���?��Qk$;GI�㋳�B(A���SQ�y^'��=��IL��I<����8P�р+��IO]yw*���W�㵦� ��ʏ|+�=�F�lL���i�v;��E�bߞك�E�w���;�;�����D��d�q�E�8� !�4�Y@j�*q���R��,o���[0��ۥnW	�w�ݥ�	�����Wr���o�~8�����`eis;]���lS�[t+bkYT��P+���w���@ ��n��cV&'���X	6@�O<%	`3��U�x�|�2k�|xFWZ3�4[cShk%綕�_�x��
B�M,&Cz.9�b[_66���O�-.�c���#+���r�n���?������������� z��~�p���M	BKil�I.��:2d�K�`ןW�m�؊��Glw�E|��*}C�:�]��>bCw�HcU�,z@�f�
���)n_���˔����5e3�Ѱ#�����ѩ���u��=sB��D����,hR��&]� N)`r�ۦy0���qG7�@�k�J��o�E����#e͢�Ong�P^?�&��)>f�Ԛ�VP���SyX����@�T�ƌ�F����܉W�Ae����A��V�2��q#�e l���}DUuh1V�_��*���L���=0�ɷ���%�I?��L�貚gO��t�<���$�����²( ��I<ϵK�dK-�o���7��al7<���~,7�9�tݖ���\lzx�����Q��9mk*�r� K~��Z����� �����_�\�X�oά�}�9��5!�ޭ,���ueU	 (T
m�Z�UΟ��,�������5P�#��T�W{'�c����\�	�Y���~������H��Hh����Hܧ����l���I��/&��UML	�����@�u�ك�j� G��Ҁ�Z-�=��]���э@���ֳ*D�A����N��#��������'���X���QԒ��o�J������ځ?Z�Ȯ�����g��Cbq���)���;c���/H��j;Ef���	r�R���Yb�&X�G��{sES�T��WX��_(@'���=�>UO؝H�2	�_����r�˰��$�\�O�}xJz>�-�5o�D��a�0[G_]W����)�QQ�U�D1t�Df;�4��,�!��v��-����j����Y�V���Y$��O��������X7e�5�=k�t"��'�x���7M	$q��۶��u�
U�^"����9Ǎ(�Y��]�x�������q�����Iʊ�?:q�Zrnm+�$��u6�r�1J����W�CE~mZz��d8ރ�V0T�v����XI��0ӳ�b�>��[;~;XUt�H��"V�a�aF�@��0%����/9���L?�D��CĠ�Ya��ڽT�w�k{T��MЌ�X�b�?9)�[s����>��,�+��[�w���ず��C�cj����˺�T���^v��Fy�H�y1K�-�����-�/�a	Ȝ�5�g�!��Y\}�׹i�|�r��FƆ"_]њ�l.�h���1I�NnD=��-�����k7�}ou���m���i#5�iZ�-S��y�2��u2p��l�I(u���:#l���k����M���n��@gP:�B���i���6�0����6+�����v�qJ�8�18k��F�󏺁��$���f^tl����%9K����,3G����W�)ǀ5�p�h�-�q�ԬWY�ut|�6pQȢ1z�C�f���S�/���c�����/��Mi[#�������f��r�� �=���ز�4��b�/����_U&�V{k���j��7V'M����;��J�2��m��k\-T�K��n]iF��I��]�Mf�gg���[�A���.
HF.�� a�!܁�����jv��a~�@X��D�MX���mBLٱ|W���>��5���ch�Q�K�ynˈ��l� �"�?�D��̮�^Q:��!����Jej��-���[$���OKI)��;�sB0��˘��nb��q������c����"�`.�0���>�A��h��7�8�U�ڞ��o�8R��٭R�؋��T��0��|�]`�ʁ�{r����9��oڵ\F/��:�
�׳3��{h�!����ZRBM �ɡ��,q|Y�d�H{���= ��)c*�
!`����E��(����r4��`��3U���sd��ԝ�Tw�LH1�Té0�$�9ћ
��"�����pl[�O�t��M�0�%LR�^g��2��6��@~�I([[)�WW{��=>msG����l��d�Z���+�=�x��Lp���U)Zմ�ؠ��H](U8y0ܥ��p�����gK��LD𺟔����j�Mٹ����B��l�&�1���w�\a<78����q���I�����@���"+�R?0����t"���,�\x]�IS�����fyV�E"���t�R)7�D?6'�R�C0��6X�1k��3W���E�ؼã5�ː���|cG/�f%jxu��Tf��I �T�R�x����tU�Ô����Y+�jw����8ߎP���՛���퍸n����#�5���Y 9c�?��v{�Ŋ�dȮertYoʼ���I:h�Q[h����&���ߍbQ����P�z�w��âl�۲��{m�/^*.\�rc� DEdAT`9Ԛ���c�4@�;^�L<�J��Qc,=����}�Y6��O)M��2H���ė� �M1�D{���T��~�p�8'�g�-{^��cҾK$��U��FY��\y`]Io9'\�� ;m�?C�ɦ?gK3R10ڣ���z>"a��O7��7ݣ��G��t�0&�RUq^ڌoss̈́�2-�GED��ݻ��c�ݛq��ԕ��w�ZU��D��h沏H��Ľ���n_l�I��0�\1�I�"��y���Yx����B�(T^s�.�Ҿ���P7݄���`��w�=�5 �3�����_4�]^�)څ��YJ��F�����p���Y援ڟuɗ���>	���l�*za=}�N��I}��_��Š=ɹ�8?�[����E��f��Ć�.Ϲ�f^b����a>��0����J-!�u�㡽�eR}�����D�,��|��	�j8�W�K&*�����XJI��r�HK�z09�G�-�:!����x���qr��te��f���RUkv��0��p��G<�Ur��j��d|�־�וl����
+N�<Zƃ;{���,'b�{���)�����/^0�&u��>ZP���Iz����љ���uY2X�"�)��8_��,��A��W0�1��h9ܻP";kq�դ���r�4�%:�	!��ؐ,r +�E�${48���.�1w:t��ə?5����d.��#u�*��a�	���s���x�E��Z�����!�<p�bi��M���R�*�=+O�'�&�q|gU�����s;����xF4��'sM�'g�!�<QSEJW�l<W%K���b�)�%ҫ��{�x"���]��^o����&j^��䶣�Q��雙͊������,��l�W�j�q"el��� �c���� �3T���{ѱ��̡Re��z����8�����Gq'0!�T����s����vP��,�o#Q"y, �0�f�V�#��}M� v��)�[����7�VB
�ڣ���NY���73֔(a���0�[�����)3�1Vۦ�(�u�EhlRc�NDx�?��A��5�)d����e�`*,L5� /�Ɇ�tY�>���t������"��]�;U�dqg�o����ݘ�G�z�z�gSL͕4�����{��$$�pyCK��B��H�'Q b���pK@��@�Q��GD�&��W�4�����w"��H���HF|���5�xv�B�I[���#.��2�LHt�M1ml|g������8,����Mv�_(d�����u�ɺ�."JK��V'ښx�� ^fe(��i�T�)��S���E����P�5�J/���m�L*?���c�֨a��I%"������0��_�k�j�Ә�Mx&)&���i�A��76���!f�th&K�"b�yYl�6ޘ��ٯ���|�Y�#��x����ȭ�|������<�������*�^���c<�	����7q�2Hn~)`J��Q2X�@i֪�,��.\�ɕ�7��XG�����kyb䃤��X��"�&�h�px<=�}Pn��=����d�c�)I��H��\�щ��ׁ7k��V���Ր(C�p
��O,U��o0X�پ4��z�q�JL�q�*'jͨ���d�`/�I=����2���)�p��k��Lr	�t��O������o��*�-$׸�+u�>Z!���{\V�3�Z�I�1P����ů'�I���AD�p�����Q������i�<�--�b��X'q����̱�o�f�������!��\�?�{��f�t뾻��T�7-��O����1�t˸�O|g��2B�	B�!�gG�R>�j5���{���~1���c�g�$����tk/�/F�#�Lf�3�{�BD���Ć�?���G?�D1���&��^�����np�Bh�,��9���ԷcS�ԛ�3��:��S5�+ERN�}]4��F ���eov<����ɓ���g&�?�"�RA���)�랶�̾�(bN ��?q��7�����`��p�5�����S2շ��+�aL���d�����~i�^l�����x��>6�稜����(�X���wJ���]1���Z][7�{m��s�f!��6pC�8�jP����k���8�?�h+{ci��I2A�����6i[�n���oW�5�nR���?S	�x��(��Yh*����Z�.���$���[ixg�ƧB�5���1��H�����f ��(�^q�z�&d��M�㐉S�Tm��W��A�L���/� '
�fx���!�=��b�`72e'�`;�.��g_H7Y��r<qOo�{�XDGg-E���w�=�Fb���a�J�]lц�\!K��a�룝�c��8���H8 ���A6;��"Z���<�q�x�#��O���Z_��6�Ҧ��ڥ@$kК=%�=�Q"A2m��A�#u����f��`�@Yb��G�E�.��pa��x��ap��J�<8���!�Ę���E#��%��-�Q�Yu���n�S�IS@Kم3�����^�1`8��ᘳ�ZX@G�ヌ����PZ�ӊ�8a��A�.x'W�m4N'^�U;�j� D�"�8���8��0�*��΃\��l���UŰm�?�Q��Z.��4�`��� [��?�������6=��U�d��X���l�`XJ�Z�'�|tǇn��]��K�IpW�L�ɯ�+! ,r���y�M�V�H+l�11��L~�InTK��Max�u��zk���Y���.|���u.�wtm��& �/�jw�����E�=s E�����\R�+^a@V�.w@���K�&H��Ȉ��� (!"w�1�s���J@�Y�+�`a)��X�����m_�?����}���H��O� �,ٴ8G&D�@�E��%A�d:�SN{7ьL����֝��NR=�<���CY枢 ;�M:����CP��u��fT�:���bJ��	e?�	��SS����[f�Z<�o�*���%��i�+�Zg1�:Ѕw�9!fe=��T�5��2�I�~(U�X��(#]��;s
_�56�)���*����z�P����EC�	��)3z���B���:K��LC`��N��k�8�?�	��g���}�Ә���u���〫
�Ԥ��I���<(���I\�A�jy��/#�;z��V�������������ٯ{�cx8=iw��~�04 aY У�2�z�j~�zEq(ƛ��1��vg��?�_����a��e�~�5+f��}�ID?��\l�F��]�%7C��ְ�	]�| �*��?�>i�ĬѦc���I���i
h=����%cD���s�wE{��hFzس���#��6O��O����u������ a���M��S��l����j{oIZ��ԡ��}��V�,# ^͊�Н�n"�$H��HV<n�������D7R�~�zn�?�R��;vQ�L�g�x��a�V�u�7��V@���6����X�>Q8VGY��=4����еQ�G���g�'E�}� ݪI���	`o}�ca��\R�Ʊ^]�Q.z�3���O�1Ö��ͺYK�N0,u�^�KZN�\ �A��{����k����D�+�GHj���p�!Z�*���z���zB!�o���#m�ܴ@+&�sރP̀&����-%%�S�|)�<\�9��������7m/`{��%�?�����x����{-�S�n�O �-jPv��]���BI[� UY0��=R�*i]6=:�������A�~�$�G�?��D䉐�1W�������`�$I^sJ=����(�u�(aJ�	2R�"��5���a1� FKb�m�GG!�/�yѦ�6�Ε�t�r�`v�z���[��)%_��p�t>��!�2�E�z�%�6D͑[K��B?��r��;	�VI�Jk�e}��ն�"Z>�8
(Q$�Jkxԥ;5Tݧu����l�t�x�:)BFR�}J�#�
�
�{T��P�n��+S��4�δ�X�����2�z�8i�*Hc�F�rS�K��I7�UT� ��hab����L����9㉹�����Dt�̣�Q��x�4����-��̠�4jٰB`4�H�+ʨ{�#��c���j���=�R���Ψrs¤K�%[���ZZ�ޟ�w+K��~��y�\�p.h��iy8���8͟��ڨ%���I�$Vh���]����O����HO�_i�f� .����ާ���?�N(V�1����C��Ί�o��kMo�X8�ψڽ��U��G0�]���ݔ����<�����;Z��c�3��,�Z!j�`K�`_�J���>Y��s��G�t�Ĵ��9�>a�B�cGz���cU:���L'���v�ަ�S�Vάޛ�0+
�����]X��n�6�J���,
�����/1Rg�v����W���?M������z_���:7�_,�j�8�m($�
`�7h�O���0۲��r�g�����e�>�.⮉_�l��J�gR�7��AĞ����f�y����<�U-������[�k`�q��_:�#���f���,��F9���d�I��o�*�6z��s�q�r��sh�E88�YB V��ò(7Ā׼i���s�=jꐹIխ��D���C7Y *�E����ұ[֬�K�+����4y���^�	)�V<M݂��iR�|bs��M��n����w�\��IB>C @�Z�8��F�P�5�v4IS>�vl�jKo��n����-�Ţdin��ke�{Ɣ�X�#��fz�ѰQ{h����b���!K����B���٘�cjh�,�'H0�G��0�u����Z���O��~��}3JX�,��I���2#f��$;�6$w��}�y�<��sO,��?M�2m9��m�#�P����n��y<�Ir�+yn�W��W�a�:�r[��e��k]��D|^�̶�A�=�}��&�;���N��omDXP�:�hx�V6X�9�:ˊ@��ui���D�l�
��1K��#$j��T%>EK���'��p�*At���n���������y%�.�g>�&6���?Τ_�J�w�~�K���ށ^ES�o�<���m�kF���s���g�Ӱ#	��_�f�
W(i	Fq!��'V@���f�yD"�^{,���x��'�/q)o��z�obIc�2s>M;��ȇJs�=�|�<�����3d��I�Љ�_l���Q_�[n�p@�T�Sl�dCsZ�A4��'l�?i�Qi\}�|oh✺:�s����	������R������w˕=����߱����:�18��j��dmnť��L7���|hF�x�`u�f�����i3��->xN��w5��^�ˬ"���Gg�+f��(g�9�ݤb���X(���v%8���?�ى�k��`⼐��y׷N�*z�2JX��B1O��T��p��}�ϴM�W��K������wd>W%=��Y^�� ��M�lg�]zy���fVn'�'���!x�*��F�(m�1���oi�e<�.�ҩ���bq�]F]� ���6g|u�E���ӓ�P���|7�<�b�;*r�p��Fd)@D �<#�Q��k��y�ݍ��HgČ�fy�� ��)>������5қ��\�w���㖟�	��w1g,�b6�?��Y��tf������4�LC�5,�3^TBw�f[٦|<�͢�8���aφH�?�7-�	�ģqxIM>>�&���'�Zb9�OT�-\H�G���o��_Yq�� 전MQ˻�e"�8�@��W�8 ש4N4�L;Ӯ�����C'|��xb���e����X��m��΁����(P/���"�X�Y
q��\a`m�o��$z4�ܥ��Xc��Pݲ;9�kw6������3�Z��AA�U������I�o�=���-B�ԒJQ���g�WE�_�S��Xt���q9��q�.���H�]�h�*�7�c��\JDֶ2�d� �y�a���2�����?W9��~k����:E6i��������N ����Q���>�u� 1��#���Q!Ԃ�YO�a����
���{a1x0����{K�"D�X�P��������o�n����YX�~'�P��΢O����)��E� c���~�(+�C�ѿt�ʋ5����lA}��i�v��K*"��*r-��=EN��N��p��|\�
;�qcr-=W������*ȍ�)����O����Gx';�|�W��duP1�^�-�8։�sΡݸ_ԑ��X`�n�x���L���3����[�Z]���`�O�������5�y9�(s1���̈̓e�>��Q�q��p��gA��%.Uf8�`۹(��ꭽ�δyc
`��_�[9�hKD�)�
t�E}���c����t�o��^O�ס1M�EC�{}#� #��)�<lz�pa��H���i������iQ}ś��ժw"���������'Zh�5��0_�E({9�F���pb!����9��~�M܈W=
��):�q^@hCzxT̥iW�g�6����� r���p�C�����7�����F��z=����M~;���� #X�����Lj�y!������gE�8�O0���v�|��%��*)�q�C�훯R��-&��\⣩���'!Ɏ~��G�`��8!��O<o�H�fA��A/u�q�DQ_�N�IO� �c,��}�"����в ㄩ#T����th*"�h��j� ���@��v��r�u��YX�����8Ls�V�q2�?8ŋ�SgM��S�U��Ũ���b�NdV1�h}2��|��9���ZҏII�����y��ᤶ[c�_]���~��sJB����E��Q&�߹�1�Gf$�i��"�Q�d·bo	�N��G��O&��N�I=��>�lgw>%cI����G� p��d�m%��������I�կ�Đr�� d7��	W^�E�~WLL2�:'䧽l2��%s.Չ1�O��y(1�����J-�r�5���r�M�ep�D�ǹ�r`4�<� �d��x�E�WȊ-	Ad�D�������
_k��5*@A���d����U3���Áh
�Y����a�nGie~6挴R^PS(S�O^bI�q��������F&��~j�^�����>��{d��T�Y��3L���i�ٕ���8�u�Է��ct���6�6�����%&��gn�΅��L��������5�-2�g��=2��$���j�����U	��=O�*h���B��ı�z�W��B�jU�0�э��`���F�l�i�~V��s�n�4�F�"gD�Y���d!�N⸇��J/7)��D��y١O�K�p�,&k����A��_��l"9�T��AA��l`*ϖXe���`�9x�x "���I�c3�!��Š���,���N���Ù �ˏ�

������u��{�g������Dp����^l�e7b� +�l^��>m��I�?��E���;O�qШ�[e
�q��>��;}a�A����&���?��ꔋ'�OiznO��;��'G'���2�2D=p9b��?*
�b8"����[�b�X��=��kI��%ԌȽ\i�UIs��b���'3P4���s�ͧ1�lI���Z~ز�le�Has�����i�,M8w�3Ř���B(u�xJ�� ���FfU=�	3�Mb!�.���N�q�A'�$d��b�1�Eщ$���h����]c6����U߻���}Yk��*>�9�Z�-q*bE��e���ew���sz�(�՚�#+Z��_�$���ScݚaWv�Р|?Z���TTq �Z�Y4�J�'Aښi�2�����(k4�<���Z}����`�$�>�_�^# ��e���#�_��ޡ��6F��=8�$s@�@�7/��%kzL�9�����.;z�Y�+փ�Fcaeg����v�aY%Z�;�pC�+��R�I�
�.��:ϳJ���H{��[�H���nK��r$%
m�)M�8r��aaSY��}�Y��	�&?��T�s��������A�S5��N�N�{�6qr�ɺ֭��pzK:�J�x�t�/K�l��gr���w�}Vv��Bv���s�I����'Of�� 2�8C����g~��+��������
=���M�8��z��s5G+�6ך�v���H��g�<����	M�w��_H�����NPi� %�k�-!<z���#f�6�Ʉ���������2�ײ��ab�N|/�[`��+�B9ſM�sX O�2~�5+��I1�cqz�[x��2��^5�hʃ9k]f��8H��ʔk2�1-E.��}޻Vip��EwK��(A���sIa�����<.X��9�MY��rn�<^~�� 9GP~�'��H�G[bKOwiL�T�˺�.ԡ�/.QJy fk�@�3���� D+*���ai2ڠ�|�N`��3P�U7�jտ���y��P�j�<�2; 	կ��\U�B��?�l����T.������ _ũ)c{�t�ʨ,�/���]}1���r
�\�L�W�p~TAѩ�'�	�7rΪS.����>�|��s�e�_X�n���1V�'	�+hHО��(Ю��z�ݜ�!Ј�@�&LȈY� *c��.	�	QM��U�����:gy�Q�����J=���;�-�ZE j(+bT���� ��l��P��	�Imܟ��H�ξ��솬�L�ˠ�"�^�h��ѨQ��Ek��O��n��r\>�
�BrAy_('�\�r�dK[F|D���� �I~�oFD�TȚ'[���b82���>���oNO�R���d��\��p�d�^���K�yx�s��nFˤ?�fX	�&��;¯�dE,D��>H�?`��+b����諢�d}�f��H�3���tɋ]zn�<FN?p(*�@��E;@�c!��CzȮhz�,P-�G'�(S1�}9�|�_s�bBug�GK��@}�����;����6��,�O].�|�D��{}�I��#��Rhz�j"�`�un��`X��r8���t�ߌ��A��bm��+�miM
yk�}�L\'l*��Z�G�9q���+,F���,�3�~%/����Dl��������Y�;K��'��] 8��"��m�~��z�B���ޛ6Pˎ4��|�^��"���[��.^�e�0���ЯwL���/����e$�
�E<LNX�υi���b��8	�p(/��uZ���a�^	��gz�9֔s�}_��y�8�m�J8��*u��ٜ��KK�|�kt� (0��0!�;�7�G��j�c�V_���󟓓
��1�������E�_��kM6a'흑�,��+ʱ�!VG���~NY��=�%TDНR_���{��(~8]��I�V AU�X�Z�x���-v_jH8{�����u�y]>���������K>�\V�4\�|��o�r�V�Pl�3Ii�R ��PRG��"~�%�~��ᗚR���J��JA ��;}�z����1Ve0�Ѩ��z��m��åL>��3��Ү�[f���G�R7��v+��KD�s�c��C����M֞�U�q��ğ���H�k��L��!������:�VTM�t�7�ٙ}�g��NJ�5���UǯF��@1�P�_"^�%Ɨ�TW=�Ӱx{cZڣ�v��>��i�j�D�c:��֙��&tPy%K�躏��ԃ�GN손�I��h�e(��!b܋
��0os���=�¥(�~�I���x����������j�4�@L��}��C���r*��j57c!;A��/2aʔ]� ���
����=6V����z)����������'W� k3h�k.�d��o���V)-u�?����A|-��z�}���M���aR�\���T�R���%������N��m�!�M9��ׯ�ȷW,�#�t�Ge�;�e��J�`v٥�Re�D���i��&~i���&58�g�n��%���^�c�+J8P.b���HY\�|dQ�8K�C�ƽIӡ�z�w�7dL؅�gqq�Q����=�̏˂D���1���-�9B��P����Շr�����JS5�N)�G3��:ՄM�*'�J?��A�݅@���5,���}�/�1��W���b#�?��f�vОy��̨���A���E��Rl�KO�O͵��^q��!����(8}���c����I}R�afD$�Iޱ���c�_m,18=ϫ�
	���\����圉���]cEF�2D�'h�h}!���Hv��p����V(P�8���L�_S���\~��o�wU1'����8���
�&���TK�;�j��rN�(�j�烆?��LBE�ƣ��t�#��wCA�_ST&�b@��jOt��A�@�n�L�P���0{w8���]��)"m's���?�A��N��:A�_�"��偡vn�e.{��4�oV1R�%��x�y5JH�a�/RI18��t�jZ�\O�A��Z�VԔ��_��~%\J��Jm~u���~��`Q�k�nO�S~˭a|Қ�FGÏ�4�iQ�7Ma��857�:9Y�R=p�}���¼}M�6[��:�E�RSyaS��y�@���CH���e�9c'��h�{� 9sD�T��.cV�V)	a�t���IS!&�8�j�"�ID�w�O8�=�%���4����n��t�E��nh����N���.v
b��z��y]�K�y��]��O=[Q�K����3Y���f����p9}y�M��$ 0(��˙B�eJ�u
f�O��������/���=<�TG�⸋;''�=�ao^������ܹWMY�G;��/ї���є�D��<TH��6�V:��G�F#���U��YK�-̗�=�pW=���J�:>X�
8002i�F �¥:�J��%��o����A̔'�a&�����F�W��Z�+%�j����
�(����pPM2V��x8&���J�!�+�u��(�ٚ���Ά�\�I�!�ַ�,�d%vHsq�f��5�e��k1b�I*u�g�HACK ����Z��Y�䰞m��fN,�B^$5O%��pj}auJ�@	��)�bi�I4�[�������"ST6ctM�β�}�'`��P����1���G��^��,|�h�9�%�7�5eA��_�j��P��T�d��O��^�������ء��Dǹ=��/�{z����6;���t��-�H3�7|AV�ˡzE�8�����'�Ӂk?S��V���;�7E\�ɾM�o��~����\��� `G�³��x��"��Ǐ�R
�-n����%�ƃ�X�c�I!,�Ŧ�=�����,k`�<V�^�$}(aSN7���b�n|�E���n1 ���<�!�4�����mFVư���mZ���P>���wAuApuI�%OLF�9�|��Hf��OS�:W�2�sE ^ˆZ��HaܜFx�^ad���b�1>ؖ�Y���ۨ�C���ѱ���>��`�
�Kǵ
�� ҁ��������+b���`v�OzB�Hv��tG�pP�xeB�m��fÍ4y	�6p�tC	�)��QL��P#O�i0��{�h�t���i��GO��ұո+��栙-��M�,o�V�n�÷�!~��WӍF���_!��4#�}BS���bGC��+0
�`��f)�ww�� qU��b�~I�d�u����).D�n��`�(�M��#�0<�*��,4��̓��f�Ky$����[(��-��pn�0�2�-\��D�Ic�#���Nėr�=k�?�D�7�FV�ޓI(�s�	�J޾�mW�~�T��xZ-��Q7a�)|���[F��p�ȑM��e	�����!o��䍚`��s��9'R-x�����;�SS�'�'�ĸ*�n�6�7|ф��r�U�yx\�r���X �c*]��d�UY��7�i�8>�&"��Z��RZ�U]��C�'���F�܁� �Qz��óm`���mgA�8!OU���	���WY�����+�AiE􌴋$�1��K�L�\H�Y��1;�������C��D�ZA��)Q����ѽ"8U�2�C���#�-K|k��ï[A�s[1�GU��Bo���hN�����U}*�W�ğx�al�[�!ʩ&�S VE��#7�q�E�&���V1�,�H
7fH��?�T��>�<���
�Ǌ�5@y��}d��p� X��b�p@+��m����� se7���I7�An6po�����K ��*��{�v�HF8]s�����	s��'�|��s�
>��-��Y������!��}�Ky��ׄ>M�;��l���L��Cn�RV�/�{|(����]6YS�[����
�p&�|Y�Zxg��J�a���*$���F)��(u�T.�$9��e{�8�Sy������[m�6�G%������e�B�o���X�v�?��!��1�׌�b-;Y`ѳqh!Av0�z]���HT�ޜ�?��t �I#TB,
����~�vi�e<U��nD٢�r;M�z�uT���=���9�NZ1�o��A��눙��[@@�XG�z�����\��{
ϰ��i�6! �����#;��%�Y�Z�����/��Ɛ�X�D�S��X�XM��'�^�vۼF�%��p��ԯ�qM+���Ky�:��k�$b���+)�L��G�an�P�6��1�������
����~ΣO�)
�"0#y��M�oT���Z��\N�cӕ���h�`$ӌ�]b'���.��ށ��b}�^�y����'���=L��_,�l_�G|:�I�R�.��(�D/�[9�ct	�|m�Q���v���?�� �D�� �����"2��/��szv����4w4y�L^L��oD��]��>��I)���I��/_�W1-.?eR1��]��IF.L&��^���8�/n}KVV��7�dv*T�n�j��lʔӂ*fT'��Pa�[�<7`fҊ�չ��6N�i���ǴÛ$T��!2��Ij4n��שEf�13�Ѩl�a�ل7����E�F��H_�71���Ɣ�=t�{JvZ<V�y���V q����5$�Q�Q��Hޜu];~g�t7 v ����PP�o�	�6��`$�%�~b�3�y��m��q����5���
��+EÎV�r�\uZ�,���Pԩah
=��U�;t�h��C
 cBE8/A�g���hu��Wf��c��$"c�r;��׉wql�^��px�Y�ʶr��lWE��l��7�6%��z�N��?��4�:�23��8�)Y����Y�Go�P��C�1u^
������	$��h�z���1�d��c�,O,��+�>��L�*��7�aP��齣sɪ�6��T+:6��D�ޭ;���$���g�}H���D$E�$�T���D��Д�q+D'�%��x�(��d�!����K�WSnqrpS��td}v����D�Yݏ�_�!v=��<���j�v�h�d�x��f�JL7?Dg�`ۺ�6�lH¢U	�bK\��c�N����ڧʖ��Z��jk��� �E���dF$Q�}�����
�T�8��R��^�Ms��ͷ},�})�&k<�㙲�u��m{�J�=#�ޢ��A����pL7�G6�4'H���I���4��W�@Rx��jj�qUF2�~�7���#Mgw3p �(��76ޚD�f��Mh56Iv4�d���q�9����ۘM���U��������23�bMS�j�u
������l׶�V�c��Kx��ќ�@�9����Y��P{ܥ�NV<��N��P e�Xm���^u�bk9P���y:��*�Qܰ��o�!m����<��@]HM +y|Ni���kM�,���O�,�J4:�cb�����mj��3��tG��Z-RI�ձufA֐X!Z�L~�y�T�?j,��{JP��Vd�R�Q��_�/fZ���I�_�Z�ehBr?��.=�,K��Ǒ�+�㸏t����0��L��a��b
X�zk��@�hߜ���W�n���F�!���Z�8��<����19eH+�{�˘�����#/��>'	�K7
uA��>�1����7�HXMե�wJ��۬����p�k]�T�/�6�r�8 8��o4�l�M��<F]����ξ���mj�T�B���R nw���;�꩟�a��˾~�������\G�ֽ��r�NN�ʊjR�\���e��J'�!����������&�p,�@����{A�>aRk#���z�YS�M��d#���`S�b�8я�V ����/.V3��ۯosԩ\���֐�
H pO(�Ɠa����Еbu�Ѡ�y����0��m�x��sQf{D�
~g{�y�X&�p��JV 缭ǁ�6������G���q�Jј�޷s"�d�ۛ�-�)ϗ��u}�-;B�g]�k��ʁk�Nc�Ul��,�m_%+}*/Be��~�Q��7jc�%a^�.�L�U8�aB�]q���z��}
	�D�l�[g���T�`<H����ȝ܍�6$p5Y�%�;�,S1�uA�PH< �˓�/��)��V�E,$��F|�Z��1��/�T  ��Vʢ.�����ކɨ�ЏI�?�u�a(3���*v/@nJ���ʂ�w��|Ǫ��Re�w0��7OHKhu�E�jg�(���-M��fv�K<.�Q?�V��A�!4;$f�|��*��ۤgM�����&�V�(#��0�,.H�!,T1��i�F��q����A4�U��޾��V5���>���K8E�@�2���Ơ�"�SU����"cU�V:^��^ �-:��,>u0������)�p�e�y@)��m�����b6x�ƴ+�⥍G�`�mFBf�@0�X���9����~;M��6�3x,_N���Q�*2^vԓIV8��
.!�Ip�D:�a��c&S��f��܈i
Qyk��m{ԙ�H�e�^^m	�����|%��Y�e���J@unH��^)fu�X��lamP�O3����ͪ��� vC1m����n����&��Q;��M_�c�B6$X�"�:4�lр�\FxΖ�E�C,|�� �1<��$QsY� 3�X�H���l��4C�>��+h8Y\υl��E�`��2��p�d��#o-����A1MF8�X�I��J���K�N���8@[נ����Zg����V7vX���q� "Oq�5��1���qO�@[�\�Z͹�&���Ji�\1�"6��<��@���x���wa��.2��ԍ|�g-�j_w����m���tp�Y�'K��|;�+w��$`��X�ns ���`�KU��e�\�6������n��s�LڢX�@퉭`��▶:�Y�!!m�ZUJ}���0M�کጓ�A��;V�#�t��p��^4��]:]Ў����7�5ۘԬ������3��b:�{c��j$o�7{�;�R���s����a_Y�
�_��| B(vI������zk�^k9I?�3�|�c>ө;����0��r�d�� `�@��6ْ���� �ŋA�6�V��h�_�.T�1�Q�/����!�zI����cړ��B�9U9]�y�Bi�' �SS�s�b��}�]�#�O�$K�M�}��[\�yIb{D���#4Q��$Uy�;����
.nf(�v�7��&�W���O]�іq�K�9�������%$`6����k7�_�V#�2�]KC\��Y�qi�`��2�x�er�245�*���<	��������O�������������T ����}V3�y������>��H�#2����hn�U�8:֤��f.��X<�ͤ�Ts���h^354 �\t��B�G�p4���K�'50ҶA�>���^��TK�h�;���Ɍ>��8����p��o,-��������G��*�����*
����&��%�� ϣC�pٝf}�!�j�p'�r&O>��}V��[m.	P��?�e9�M1���Y�i���"-��B,KG(8���Sbet3��a���@�("�d�D��1@j�v-^�+�peq�%s����m�@�� o����Z-�^��1�k]�E�	���`d4���Ǣ ����(���n��2��
��ݴ�d�7#������;��0o}x�$�����r=�#t��@�����m�xy�q��E	�XԢ�2�6��nz���*��HpzI��;�*�l��ª�}��Zci�#C��M����������m�
q�bBe�~4�ەo'�'W�i���"���(�-�|�}L`�o)���(�e�y*r�o2�:�]��\�m%+q����@�x�G1]Ġa���?V���kIӁ��ѵ+�	��^�3�+6���E��i���[m�}��'���iY�@�o4/�)x��S(d[Vk`�j]1����X5�������ʈ�v���J^��e#�%�1)�&�'S��E<�� ��q�&~˔z�h�q��;�w����WGG���U�K�Hٔ��
���l�� ����s!�M�eZ�X^2��6�y7�k��x[�Sq�?H��z�o)��!v��V��C'M��t���k���Z�ҝW�lm-To��͠�rA��l���)r�0�O�˄�=��L���y[*b�!9UڊN�����5�r"8iS��e���,�2�ò��&p��K�W@�!@
z(�\hdGM�+�ER��D^	O/�/^{Ty��c���*F���$��ҿJ�+�_Z�K��S��~�
 �G|�_�>Ia�o��nN��%�� ���c�'�N��n��-�鋷,�O��,)8�$��{`¹�a2��!�����}�eg�W2�z"3��+*Ny@0�d�p�e4I�:����i�x�����[X�s,d���C5i�Q�23uh>%�<��~ ��X�|�CW������x�A�dw�;�ҟ�+#�O�{�_���2���������ir���䓇��,��,���WokT,��y0�6��~>��47�xj>c��4a��i���w�����ߌ���(	vd�j��ۘof#���qt�Rx�b�\�7�������?�sh����II@O���l�%��n����)8(�?T��R^�=<����^�q�n���&!{�������Mخ�I�>g� �yP�o�շN�4��"��Hm֠?!��27��1�INhr���SǃoS���9)�V�kd��kQ�o��/�u��} X):[!(qO=�{���b�MP&��b��b=�=���b|��w���<}U�q��z�87�PAhouۋ=l?��5$�B�ZuZ��z��"}-�A1���IɁQ_p���HZ���ڈ��nY�M��m���)݈����]�M\��j~J�?�6uE���
��Z������g� %}��}HLCW�(�4�uK��m�ҿ-X�^���H����0u@"F`C��/�_�9�Q��q�(����F�]=��'���&����6i��}�-�(\��q\Ow�j�9!�����酼��uĈ�	��	lR(�IF� �Z`�agڶ��%�q[�p#Z��n�hܲ�1�&<a^q$�s2S�:u��*�4*ԛc�B�^A]�=�/ğ(��ꀉJN���$��U/Kå�#b��!$5���j����'8�ޟ�1����;�A&��z7��O�`'��a�#���1����X
ơe���އ�o�S�މS2]���j����km���0������}�T�v�،�@Ȫ�>:{�������"/	Y��4�~��mj��s���
`�t���ĖWX��G1z߼��Pɶ3	��=T����,v �5t.n��kѤ�C��矦ĥ��V}�U{4�Qk�l��(�@F�ݹ�E�e�#/=l�ru���d7ze#^S"�0_s��ud4/�C�?�����1��(f-p�.!^����Ʃ�V������(�@�s���]�$V��o�F��C��}�S�`O��F/���w�z���PJo��/� ��2̆\m/2�f`�[�#���%��`LȪ�_{�%��X�^�{;�0�lb�I��5.��6�7f䁜v)JJ���K-��{<A?�K�8sݻB�#�LBD�V�����S� �b��^ �!�v�iE6g�������?ە�o-� m|N��?�m)��,�J�+M��5�HĚ驚%�-2#� ���楻��3JH���K1}��7�����Fa�
�p�#A��&m��Ì����/5B �M��	��]Ǜ��$��5J�u�>v L��6�-K��N/a�S�1u���wq�ǐ�q���'�ǳD�
��P�З��
��N�x�?a� E�rD8� {��ʸ����r��,�L�^!qH	�=۹��mc���~����is�NˎܬCT�<-y����/P��ɡX�]�jD0���0ؔrs֧U�ڍL��I|����xv�kEg�F��΅(�����W������Jp�Rޅ2�r�$�n������k�#s�=�O�q�gL�_h��0�2��5� �T���r�:���������M��V�^PA9�;�qqt�'�9���ֹ�V�x+z<���s(ﳛ�,yF�8aօ�1���D_hXD$�*