��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&r�F���oh��7�K=]ꎁCa-\�م��p�232S���sU�4lf}�_Z�k'�UF6P�Yv��OGp���LQ�����&�t��'����>R�5P�7���h`��^�ViOVKOnQ�E�K" ��+Tn��BS�c�T�A���&���UM7��^O�j3�pt�Lq+�F4f}�n
�[gi�	=�<�?�M�J�̂�L�$0Q�n�,�o[���p�D�D`l��  Ū��ˬ��qEqՖ a�SS噯O݈��PKdAD.'�9�!Dϫ��߱����p�s��� |���M{G���S�1Z��7X��YHF#�h&��!
����ҫ��>����*p~���,f����S�U��فh+P\�յ�4"A�d��h�)'��t2OD i�)$�
����ti�u%@� ��=o���i�v�OT(�����:���8��O���]w�*��S�|�as~.�C�K�a&&b��д�&K6�GV�Zv��+v��Ӵ��pm�F�d�"Ԍ�b�m�K��I��������B�r��N���7��wC�\O���=�KXF��vcH�#3v6Q%X2W��F/�����U}a���dP��/��v�a�Ő맛�A�^�4	�5���i����z��'��Z�j7=�qGlS0:yv �ܫdUO+�+�Cц��b�1%�h7)�z��ܿ\�� k�����PN�O��HKl"��BO���y��|�wi_��]3X�˱SZ��2"	$;�(�b�2%٣��:]�%)U�	��I�z�����S>�gՓ
��y�+�O�o������U�ӌ:c'���m�v��+Ck��O�Ѧ޻]��ӾV߂�١�s7��F�)vi�� 	1���q#O=�:!��UF^�e .�2$7rz��(KA�`�ON���pƍGo6:Q�O�/v��֛��[�5	1=��Q��^P̶���}Q�D)���%.|�;�4J�����K�:%��$���>�I����ȣ���{��]� 8�"M���д*[�=�v]�`i�X��y���|���}dԥهt2������f���ܣ~_2��V�B�/��Kq�3�]�yU�TI^��^�9�W���ݎ�XY:�<�qwR�F���e�ͥd�n/!p��s��aʑ��� ����h>�w��z����d��C�6U��\rRM#"�+�AmQ��&\`�ic���O�J|d�C8��5�r�}��@�A8�4��\���V�c����*l~� :���I[bx�ǟ��ߒb
�GCӵo@891ې��8�l4E�+ۭ����#n�̈́}�� p(��	��E�z4�M��y.�*�#��J�)yt91$�S�"��a's�?j>Z�T������[2Z�FL�n�6��o���"�'������j�*�JR�L~�hW�ָ^��h�x����yQ8GH��_��I/[V,����Mᒗ���wG��i���C�]�|Ű��T��t�U���R����E� �>�y�ƭ;��Ú�?}{�d�_�����:8�!�d�� �ýP6!q�cv͂WX��Y�@�#ae|�5=�A�`tRmI7����X��tvr��r��%Z�]ٌu�u�s�@��B�TgԬn�U˚�Z�d	sn�oZqR�����/U�iZЗ��8Qn��?"������5��eʔ9"�WJ�Ė�[����8�?�"����������� �߶C^�$F2�Z��a)�y5�p�@
��/��s@��c侞m����ES�����,.9�wl%��A��Qc���� ���t%K���n�,���SM�w0tҝ�;u�2�}�����[��#��b�ZK����#��+4 �4���Ǘ���𱸛 󷦗U���_��r5굂s��D"DꙞ�pt�{M�WzpR��*jw�X�閉wG���M'����X?�\�us�����!���(iO���"�?�X�98x���z=E�w�E�/+.��[�W��r>�����ɟ�@��y�(tY)���cA�N�&���d��fM���5x��p�	����r̈�*��0���l���?ǰ�L��a�pR�Kr���ޗ)cF� �T���^���2��4���sv輆��K׻ޠ�ߖ)���G�U'~�����"sm�*!����5\�4H��r��K����O�7A�1�S!�҅��㘿��	�E6�K^��{�n�2�C�-�j�K�I��l#�ŰZ6Pb'yL �С+*�Y�J�c������]�I$���>�?�qocF���W�;h��G'I����O;�w֚Os��x�O��vJ��^��DȲj3db�Q?Ita��~�h��Y±T�o��3�N:��Z=.7��P%��rf^�ciH�;�q���;�T	��F��\�D��ف4~F\�#N�6>Q9��ஐ�@�俘��V���� �]���g-46�X�!e7����u��a�q��]�h?*�7���֒� ;o�Z�4��*����T�F�55��ht���`�F�ܒ�#�Ye%��	��oF
"�*ވk<�7�H�_y�D�|]ur��2�~�f!�#�	<JKz�K>~U�8��I��'�hf��V�`�P��3���0�N�k�@}���xJ1}�9#�N�k:�nr����D�3��d�˵p��!�qxڄސ��`�>��P�������ƀ G�^Zۀ��&C�F�K�F��6휥\ Җ�+NE��s��DZ%�3�~R��+���#�w�Y4�@gm���/3�3���d�a��q��j����!��E�_Y������g�����݌���