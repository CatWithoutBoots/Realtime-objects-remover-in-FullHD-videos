��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�Pk���<�T2���݉�a��<�B�t�7$@�}��K#L!9p��ud��^ڵ�@j��Ff{�緄��@~�z���G*FIC�����J�S0��
j�xp�M�,���*����,e�uiхq�ߛົB����>26��2J<����9V��¦�x��:� �5��˳Y'`t��5s�����}��B{��J�B��&s���.�2Q:�a�����!�2mjC[]���⊀�������c[w�M2�����Í
'~��� Z�ӵ�<'?��R`6ݜ��(I!�Gҝ����D�
�����M�d�G�!�����"�M�e��ώS�W:���K����l��q�?�s���G��#!Z4�lȿ*#o�`��o�I�

]�����)����Q��shV@��3�֢Ծ�����`S8��r��H{zĚ�ﳢ�.�TC�}��$w�H�����[�*��؉	^.��{�d�*�݈����I�4=�,g+��k}�B%�����
�4���*�\���Q��c0 ��3�*��	���F��*��߆��?�4�D2��p>���F�����:�#�D��v�/lr�����K̟˟�#;�?@���K$3E2�l(,��\��5�hl�;�;�\`�g�ġ>K;�h���~�~~AN�Q�����,	V�� r�xz�˒�h����m��
4�4 J>uA7�P��=��?�uպ�F >e�p�n7%�L��
d�����gN���=����9���2��D�t�rCZJ�j	�|�aQ�<�y�O
(]�iћȹ,��[�I#�vd�6o$k��3�6�!ɕ$'�o�V�`�R76�����$��@�k�����r�� �I��G�~Y]ȯ�J���o�r[�] ��29ݣ���n6����lSeUd�Ժ����{����w�K�k�N�8G�Jh|��d�Ō � jP
�3�*Z)��:���翤����$9\U}Z!���M����Y�j��Ω�{o}���3�W�3��U����%a�
I(Ձ`��MB����/S9�ڕv��j�s�t�EFԪTGA�V�b|�*�Q �j�nj�r��|N ��,R�4l�%e������,;��V�1���MZ��m�	�;��'�F�C�:=|<qmq�)�}�+�*�t�Tb�x���/�~.��6��� 0kr�?�8Ek��3��kL�&��l�c�	��y��x�.;}���6t�4�i��̴��f����d�e�4]�]/C�>v$7�f��Kw�ĩ9ëz�'*���ۛ��{���f;��N�~,��Xx$��u�z�N��bv0-
�"%�xǖ���Iۇ�����݄,g��nl�=4Xc�����&0A3T"qAnZ_�3%-+]�8�-�d�8����i(�\�s��� �!� /{Z. O��(�J�s�I� 'qe�x3�E']�(�q�C��^S'��F-�r!w��?�R�D�3��9�!��=K�M���=���<��������X�t�?�>��;�pt-[�$���9�]�*�>;�Yu}v�������u,��sR;���\|:�F��M��o��r�$�F"�f����}����@Qspk�����+��3�f�u�h-�Z���k�{k���(��q�	?�Ҝ��πI�K
�����~Y������	��\K����Ѥ�dȅ�io6������I�9��
��[�=�*֌,T~S���f�y�~��v|A���k�'��t�� �N�h�S;�y��c։��B7-���
�p3��L�;�O�i�gT��]5ݗc��.GX�o��"l�HW3l��-�T�A�-5�Y	n�
�mi�|�dxϽ���/��t������#��谜�z���A�ϟ#�L���.���to��Qe�AM�����S��%�]z�ؐx���Ep{C�����:�gBwv�Ƹ	rjAe������m���P��RY�L~]x�
�,�Dq�,q �o�G�u����9`4�`N�c뇩��ڛS��%�[&�Ӹ�#1fx��2�cH�$#(�TM9�"�ꟾ$]".ُ�L���vrq�DRE>�۴��5v��/H����&�����O-�i:[ �27h<��=���YԔ$e߉�Ƭ�	��J��bP\AP�,�r"Bd�ܔmR�����vh�W&��|"�i�95�e��v`>���nM����e)N/��v� HxK�[�k!�e�{�D�]�%�Zm��M��r�!���i��A��;�d�I��J�q8���B����2^���_~�r"��f���o�Ų7�+lT�h���	����bo]_��y[h�(g�īJ0;e��������9��>3���F}�<}�Ю{���k���d04V��/�q@O����n�i��$JY�
W{Zۛ�*.�3 @�6 gՎCU���$�/�z?_���7��~�W�9��8�Q�^��$DT��P�+md9Y-]Qn�fQ�q����:d���!��<uۤ�^�?�-d>��-���f95u��������=]5��X%iÚS>=�*�����-aj.ɣ��#^�Itgm�c�:�ޕ��.EH��9�Q���F�B�s-�J<����Q���{%������~�����~�'���J _B#���@��_'��#i/��ؾ��dÝP��3T���qI���h���Glwsl�%� �xϔ�d�2V����I�I+,�cj������[5s��<"f�qKu�+�)�����x
���%�A�5-�.|v��~^�,���R�!қ³�Ƹ�N����w�F�b!I��	��Q5���(-��,���S�Z��P�	kO�"�����}s�C�0,EA��c=D�E��������_�����:�Ϯ��(�8���ŭ��R-Z5c�8�)P~�|z�o�BL�~�d�h4��z�����.�!�F �S����
na����hzm����2��F)���]�@�V��T�-�t��@��u���g���U��z}�P�]�V�t��,�o3Ĵ_�����	�\�j���z�~�s#��(SPg���!3�9]uH�i�n��Uh�@;S"2��|Eyu���c�ˀ����'�QY��B��i�����|2N��5���*��1/`��-l	�zl�H��p�\��X��_����*^�
�@;�-.�nq1�rh׿��H���BA�y2���E�vv:}�f��)x��C�`F�M�h�R��5���ν|�����VMfR?���qU:[���uN*rC����)���3�sd9��V\�\�۹��W`�@+�8��{��W���l�c$Z�iFk���X� ��1Ϩ�pu7�\����"燗���mDҧ���f6a����Qnh��
�6�����0m;��A`�X�N�A�k����S3h�i��`�׌_�7���9�{a�����@�a:dxF��	�%�@��=�`= �b���7y��m��z�;0 ��COy�VI5L��Q>��F�p�{��J���I_�S�=b�y��>�I�o@i��������KM<�uZ�r?D[x��@�t�!>��8�a��
�����M��'�K�#�C�v�-%x�j*EW��r�$�K�3[�L��k��_��I[k<�����r���/Ծ}wߙ���!Y�jڃG�RLe��@�Z�Ș�g���[�XG7� �hE�3�z���Y3�/T�<'%k����T-c`��cxǣ��ޞi������d������._3���<>�4q��P�>6��r"O+t��X����yo��q�V-�GȨ!mA��}DUP�xʴx�f�IU1
i?���tM��O\�<i�,U����M�?[�c|e���5r��dccZs=GQ��uSMn�Ҹ&�-M(�p:����F�]t�k�������.��U^ ���E]��Յ-_=XFr_��HZ������?��hwB��Q��.3�&/� ׶k T����D�$(���B��1�H[Mn%Hf�aw�ʢ���� ʬ��䩚�0�!�������-�x0&/�\�9�NU*3��d	��]E�,�}r��)lO��%h7��J���v�"���;0]�M��7@��A
��Y��9o%�<�+/��������j��gv�>}�2� ��>�,���ṉ��!>d0YEB���L�Y�<�3HZ�0D����y3e��7|�7GLs��	��K1��Uo�iWu=�΄�-[eTQ���5c^��M��	%��C�JO��/����{O�~������"� ��7X�>�h�F���ҕg�*�V�R�%B�b��
�ʏ�Ɨ�(dɎ�Q�?�~(Y�E;�P���5u����pQ����(�#�)�ѝ�*��ᥑ�M�݅M�J$�TA&�/�6� �����������VW�l��h������������:P��ڔ��{A��/����IN�?r�9?��f�LH�о􁃭y�Us���O_IE �t�C|����CT�rS����M�'*g;�&���Y*�K�S��r��LʱK�%w�Y���;�a��O u�A�2QQ�ۡ����g	���;o�kO���� x�A�zO�P?�+�.��s9����G���=�!킴��Þk�����f/u'�m��r�y�
u���4�"�K�Qk)�a���ZF\l��A��E�����AP��lEʏc6�=$?S=���l������5n^P�2VʱNJ�Xz���-���,�r:����!�����CZ��0�T,OV�=vA�x��^�B��3N��h��Z��`K�9X�@@C�9{H�a��r�k6k:�)i�2^�N��He�́qQr�8���u8)S%bFN�eh�ij�ګ�����Zb�n�ZΊk�ǅ���j�s�������܎ݍ~�T�$�q��C�z�<�D8i��HV�tYaE�7�ٙ�ôyZ�������)r��#�U�_���e��_�^D5˳�zA��h�9�G^nʕGȢ�3a���
� �ꄎk�(����0�s�.��ik�A��dV�-�2�$(�1u�O��0%:RTCJ'����V�wel��f�&���g�Δ�f4����d��WQ�װf�&*�?�,��vp�+T-Z��E�eH��k�F5E��R��a��qoo9��_��@\���v��I7
w
t�i9R��"�2��$�?��M��Ig��f|y��*� ��(�얰zZ[�����38��݅��g�g:� ���������PB�EopS���d�������"���ne�o�^ʑ9�l��5�+sW���l5nI���zlJTpR��;:�̺yh*�"%1�'͗�=0�4b/7�OM���m���s2D����a�g�t���5���X0� ���Z��s� f��������^�2��x�pzJ�W�z�+PxNʢ�����ohVEH;5Y��j3qY�7���c�H��i+�]��x�_UZܧ�+�U����c����A��Er�'�vaK4�B�^�����Pb8K�xn�˯|F�L͒O�ͱ��YƬm��*Vp`�6� Ռr_(y�����<�"RM"ލ��JTX��n��VŊ�G`+jK��2���ց:M'�'���]���n\�MD�sO��+Zsg��qn�L@k���6?�{�U}�`��ͽ��=�J�42���;:Z?fL�5`>�Ϡ1{g�1+C�Jݭ2u��� �P�!ke�]T�%R��)�5�4~Cz8���E��۫�%���n�;�+9�����Az�Ty%ByfQ��+�������a�V4�Z�x�������	'�
�juwT����t�`X��mF&�{�o�O|ٵ���
�W��/'×����[X��rU���zdi10%�d��UCG����B���ع�W9$ud���$��G�>��_��}�f��������Ќ�>"�
�aa/i�0g����O7�2Y���w��{,J�1Xv�K�h=q���ho�!�@�I�@�Q������W��������U�I��79�����TY�T����t�Rx�d�i�˾�g�F���z�½v��H\��
�^��x�Πi�CP����̀���(T���l�4�a8+�E��]�p�`��2ڛn+�2�$(#��
fO�S��5���Cy�>���t��+��e�'=�9�t*��)����\r�j8��ٿk
\�����1d��.W�=g��'t�*t۽���ͺ%%@���L�=��G�]���3�z�~�d�
��$��ϋ�5ݐ2��%�s;b��B���5B?��c����C�`�ե��ޙ�ݔ�>���j�࿳���0� MƉ�$л��4�C��O�)Mt�|"2{r�,�~��)�����t]�B����9h�!?5�YBUH�M��wԶ�q�Ɏ��T��:�8	0���U�o��+��^1�wnQ�4"-<�� I�����{�\�7� ��C����Vԭ�cOxn
3�p�Jf_�,J��Mx��G�����x���t%$�QޱJP1�~����)e��\�����a�I���?gF&q~4Z+�3�)}����9~ɫf�M�i���'��qT��y��k-�#(F������%�Cli�c�/�mB�	�#��o��O���ȯ^	1���){*�f��#�yz����v��Ǵw~���o�u�a0~�N���A���	mJ��n�l�f��Q�������"S l���r9G*l��Gp<u
�HY����wI̲��]��4F)�o_�I�ţS�C&��"*Dp�oL�-�ǘ��D�v�ǋ�U�]�,�,�&���j'�p��}�V�}ֺ&���d�?��������7�6���O�^�B�?���q��?�ΥA�?m۫��S[�DY�j�P�N�Es���guJ������i��q� �׸{�%e[��	R#��D+��=�Gikw�4��{���X�4�D�)���W���\+�MX����A&�D��T5�s�����6��.�x� *c'%r�Fr�jB�� AZ*�Ǫ!ݜ�t�.���x`���S�z��x�V#�>
ͮ�*�E��G��mӇGJ�K�*�!��^C�?,�(�}Z�E/�*[��EQ.j���b�5e ŷ-a? �����mb�ώ"����F�~�*�����b%lQ�r���*hOE�iʟ�'������Q��J�F�閝���M�F���s�\����Z�-b�%�j��RJ'�؀�.J��Ć��Gy��:^�Δ�e��g�h�
��H�40E�6�	�ye��K>�ЄT&j쥰|�*�$��9n9S+l�t���>vP|���@�	8�1��f�i�>؆�#7OE�vL��#Ӵv��$��$x�/��F�{Ղ����-8=ɏ	�<�W�&Lюdƃ902�wd@�޷�3�w�B���Yo�k�o~=v�%������P9\�����t���5pH�#g��K?�D|?���_T���y�ԭZ��B����S�������'g$�N���rg��I�lik:ط�*+;�Y!g�tQ+KQ)vt\:̕r�zW �L�Xv�����!����GcR�a-~ַ!c�Z⬦���y���]���^4�ꈉ�S���+���B�إ�S�f�)(wGٖ�z$����p9b}B�f0Ħ�q;MC
h�;LR�jXP�����~:��4tb�s}�ug�<�]���|�a��v�MaU�j	�����E�$�l�ҘxpE7�vȚ�H���S�C#Wm�lB�+;����n YO�ܯA�MF�J����0�O�j~�e��,���5��aM��|6N'�56�x��_�4Z"� �4󥬼�?v��Z�=�y �Z㥿I�`d}�!`��2oր����C��/�S)&".V��OBT>�t��#X�?{n�)�x��1M.�O7E�
y_fV�K	�E�\4��r/��{�@��c�_h�u�l}ng�8ƶ���)��8��nY����\���*�r)^ʐ-EKA�ob@p8@�ej�Bۀ^��o��T�~x�@��O�N���Ȩ^����Ni�R2�E�kL��$��
�k/�1��/H&/}t�5lIA�$���;�u~��}�� ����򼡤���)�z�P���$3�t������k}�AT��c��h�������/��po����=(�6Ӧ���\M���3��j�<�GQ��.��)|p�F�f�Je�7�e�l���oF�yV��SM������~�<���K�V� UR���[�����v������hkA#�q5���G�X���+�4���|�{*��7?)2�AX����kq	2�Y�����;�O6�����h
w�ǟ=�/����� �t'�b1���$+&���Pb��(Ƹld��Jwh*��k�o��̜rSon�>�r� �*t�·Ѝ0�@�
�7C�jJ,�V>��\���Nt4� ^�t/�-�z/(v��oͽ���P�v�3�A�[���y�60��~�eWl��u�3�i^A�K�Ղ�9�C��8�k�i�6K�y�uI��)��+ג#PA9=N�f��/��?���(˚���\���n�f#�gP�H3=�Y{��zg�d8�VG�ٙ�?��M�r�O��`̲�NS�֖��+gf}ъ0I,1�����sl�ˎ�b+=O�G��q@� �|,d���u����{�<l��,�Fz/jP����D����I�&��m�l&�n� E�]����BՃ��R���~C{J�T�)L���G��g�ŋ�')�D�=�*��{j�ے�}�̍'��E��	[����ݘ�!t�bq1U�˰�}-��s�"i�	���]���T�G~M���fsEf
EՀG �3ѹ�q�u�]����\M�]6���@�y-��)<F	�<�}	ń�һs�T���Cf�P\��v��o~�/�������X}�$�O�FrG�b �|���O�\����?�ҵ����P�ء�2�_�V���5�/C��*�$Ц�n� 	t�����[|��k�=��X�v�7q�ݍ��$h^��*,��	B��/BH�����A�bc�O����%�l՘�l|w�j;��ܶ.�p��Ğ[h���vt�Y�=��%�~⾴���,�mF��,��7�y"�3��(����}L]�~���(@"H��mƘ��A���e�q�㭝��6I����\Y>HR;��Kz-�w ��ʀ��8����a�z�E��ȝ���;r�_��x��>!�;k��o$6�im�bq�OT�~E9�9��`G}�Yu�N&%�VɎ��'�Uά/�������B��X'�)�hi��,�,�������ȵlPFȍ��'�8��4m'�|>����'��n�lbif�P|��#�2��(4��:Q�US$��tʛK^(��y�"���� ��S��Ұ�E5�g�P�h�װ�h�s����Q> y�4�q״a�O����k"�Mº|cW��o ��j������_�yAͣH뛇���*?�,E:?)5��=�tk�3��V��^����ײ���Mj�wѺ����!���1�I"�d�*ӄ z���a��2�UE��59�Ua"=vN��FV;���ȩx�B\�Lx2���P�?v�ᦋ�*z�t�)n�5E��Q:�u�`T 5+E���+��~3���b�/,6���$���-nGvA|��Z[���rA�IƠI�����TfǏ�MC��Ju��&��@͖ر����f�E;���$TN�Ň[]u���l�eF��2�T���Iey'd\S�ڕ����V��Mw"щfG|(��p&d�v`�:���j�OB�̳]�*�����+m�~��4~z��BqpG:]����໰��`�m��f4j�᭽h��U�؈KV�
� #5��(A�T�<��W�ؤh���,�#�_ڻ/�{����9j���v�Cq�z>��Qf�ǅ�Rc`�0i��9kBk��x��g���;��0�L��t�4�SOϼUw!��'�x�R)���ާ�z���*3B��AB�Zǖ���ˁ+����Q^�P�F�>�'�Nݱ����Oz�yH��1'�:�ٶH|4�`:���H7pG5U�.�MlT$�=�0$�?zi4����S;��.t�E��a�+��-~�j�AS�K]�`���ɷ�H�{`NU(� �sݖl6�砞[�҅����f}UD單@��lT���e��*��\���\s�s�
 F��I翪4���A	�@��9T93��o<.#��h�HZq;���r�Ȩ1��G��#c�����aK�(7z>���;�����J���`u�(Ȁ4��pl�C��cNh�bɪeE)<�Ţ��	�~.��n5�u �����CZ.�X���c�G��,8ʀ螧JҾÙz�5�̒���rKW�_�M�e79���D�O�����r!q2<@MJ10m��~#$�����pm4���+B��&�1ݯ��9�6�W�����"\��S�b���4�~��O��U��&X�N�F�{����+[㬈.@��7WƲ{P�̕�AUoΰ1�ƈ
�VV3ͧ�rئ�e��(��x��
D�/����S_��|��U��3��}{�;��R�+I�R��dP�Aû�0�_��w����ͩ���Z��2,{�g�՚�B��x�Ǽ�y��s,��7Z��J�x�l*��wYh}a{9�)��;RXG@�5s됭��CX'̺�%V8�R��Զ|:��%?���wU �����^~c��y^^i��'n����º��>0zb�rj�gc��L�y��,�Qwń�*�}��[�%��:W��n��I�(�	C�2�/��M9:�/��wh�M�3���֫����X��p _�Y�7��w_;����q�)p�۳��f�˺�ȲU0��CP�k�eR�<�V��k�Y�h���
��_쿯��t����4�k%��,�h#��[�y�Gs��.�t!G�V2@��W�{�[ۨ���8O��k��]uI5m�������yb�-I353S6Ɉ�G��C�l�Dj��馋�Jx�Բ�z_g�ʏ�K��f�����db+�hJ#��:y�;;����Q�
ֽ����>�F�������s6��	+�P�c�&0���������S^ �bŦP5��CT� Ĺ�N�4/V��|ie�m@z���]#��y�X���-Z.��J��a|�y���2©�{�
3�8��ܝ���q�Ú�e�Qd7|7GI�Δr#�B8��s�/Kx������VB���5�Y���g��Se�+�|�P�R�Qf���?
�Iv�T�|���U�g��).L���������X���Eh��H�m͈��~s������Xoo�3j�������rh�T�*8�I�6ԕ`�Ī�H���&�A{�%�\wm��I��W�&�Mz�(�,>�` ��w�:MF\`�[�˭W�FƢ�z�s���|�J����|q�e!YJc��0܈��汁�>a�w��0���TMc��{�8=2]1a)!�7�b���TC4�W�-�����_� �Niۜ�n��7���oȘ@����������)m\�drd�p�i���)(�AA�H��CrS}ʊ�tUN?r=bs���� \��c�ͨH�L���|�oK�oY��75O��۞��d����ˏN�)� �~4y���),�#�V�B�cG����fu�վ��a'%�����F�\&��ԝBJI�T�x�V�#޻��p��;���-b��QE��T�l9�C��Q�T?�G���T��}�i�|>��z�*��Ɖ���"�M��:� Z�,�d�XscA��VC �1�"x��󓊤=��B6u.��ln�����yVI�Z�)����|��W�k��6����G<y���f�
-ZA~�*֩�d�,=Ru�t�|k&f����3'�U�4��gd�D�������s7w1N��˦<��k�0Ĥ��]05�FW���GdB�L�R50H�Z2�ҥ�U�Ɣ�����}����$TW
ab!f���]�]��G`�O�iX�;�U�ElQ���,ʏғ���ۇc��i"@��tj��9E3��^R�������Y:�a g\��� ��T&lgjL&4Rl�c����,v�2� ��dF���V��;�%�<]a��bК��t�QhT4��������pl�s<c�ߎ�y3�x��V�*`J���ʼ5�p��c����h��H��;�Z���c��d5X�3�q'i�X,�5`VDШ*2X����/�2��>�xH�=^g�/�w9�&r����\|�T2H�,��i�7`���䁋�~���(�f�|@�b���a�$BF�ú�DM�-���hrɏxT.	+%��ƹ'�g��;:�Oa�'�� ��q�/#};'$4�_GT�w8���Ept"~T��S�IMs�AE�098��놫�2�Y�.��hX�E�J��U���h�g��t�5�&��w)i��͖(��EBlwO�5��Q�Ax��o�tO�Im������sA�wȼ�"��9��3t�T����E~��Y����}�O���jy:@�^ ����5"�U��hA+�$G]�[�n8�,wy$�p��g��#��E������V�U�����2�r�K����Y�PM���\�Apǟ�Y��Z�&���Ŋ8`W��p���ȁ>O��{��,*�
=�*��m�b�H�ӷ��J�n^���h-#���g!u���YH�e�r�u���n�,���
AL���RLJ����֙`ҋ���1�+�7�q�\\^�k�y�D�=&��CW�Ua�Ɋ�{���*W�()�,luq�Ԑ"t����=���0�� ^�$���CX@�
M[�����C��\��^%���=k��"����e��[��5��~:n����UH*�{�x��R����9�L�a�(���T��B
��96��������?4�Mw*�7�E���i��i���,TpqЇ�� j��L����� �].<������K�R��0%j���E�Q�C�F����R�K�}�G��||������E	bӳ�n�Ӽ8����3$���:m��	��h�OQ�Y>Q������S4�%�s�G�Ȏ듑L��J�>�f(֥����+�k񞹅Q��� ���=��4�xuϮ�s��?}�2r|{��2H�� T�� 6�$g�>[�-�P����ī���ÞD�������j�B;B7L7��}�J�"�`����	j'�����~�ɍY=#���'ޗQ�)���&��Y���&��,��t1�"���'ö�?��= Δ�F�j2?b��,z�X:�6����k���&��oQh5�q�1'��,���RU5�5�wtJǯ?5�A���x�k�f�{TEt�<S�ȗ�T�6J-ɬFٺ(��Όs(��a�5K����ޝ��%��\XG!ܬ#m��L|����ĕϊi�d$�n�3�1d��q�=e�/e����r
��N�45�W��`(�-_���s�������U�m�5|��CQ#��j�Q+��1/ߘ���T!" �ovnJ�2W�wp�@�FU����L,s�
d9S�O0\`�4��z�n�P�A �g�c'�|A�]o���x����o�gt��^����C�2J碅���6�+����o�(��5���Nr^��t��V�V�g�e> �%�+@/�����:�}�۞�1W�0�M�i�y�̌	��DG�$�"�d]�����j�B__S1d�<��M�K�{���.|~.�������Q���(n�E�(> M�1��1�`��i��&`�%���Wl�/0�B,>�����?B~|�����d~��OY�.z ���4���x)"% ��[�P���`�::US�S{.�՚����Rd𫅪�( .ě�o�
�%> �<C]<`t�x�%%w�Б�bJ��S��NL_.�����P����<�?�i�S���/?�c��'Oމ�,�)��"�X�ifI �V��w��,Ã:b�А��1\�k2�lcl��?�z�Ӌ��a^�0�dK����Ӄ@&�P�,�� ��	�!��{R�M��G��!��qՇ��i��U��.�v:��\n���W�rY�G�YV�	��豯KѤ�p7|�[i5���S���������c�&�rO��f�$��`.�jh�p�xnw���T���,��k1��o�k�����ͭ�n��N�ثR�!�� ���gV�GU�����O���}F�⇫��;����P�i`���e��w�qP2ʄϿ[��!�d�.n
J��M��RF��Qb��Gt��(��<���]�FwH�:�J��1�@�� �F���p3�P�ج�a���7HB�5�v$#ȁe��C�&��B��6��ej'�cԱ�����f�#��)^��ձNaO�e���t������#���Cݮ��%᫼�2՟S$�i�1{{�)�K���tA�ͺ�s�#ol	�?n����*�u0]AFf�S;��r��ʂzsc8�����S���jg���pW|���8R��d�KP4`�կ��l�v���>Eu���������9���h�ӶH)�di=�q�+�����Q�ɺ�=�ʡoEr��ط�\�`K��z�J3�}�	k���e;%8�8֍���ޫ�HI��jx�\p��;� ә
pΗ��!VLUE>�o�I�<�0{��E�����6������A@��~����_�!ysW�]�k��9 6��sG��<� H�5=v7)�̤��R��/1}�6�6��14R3���z�`+Ć@�tw8�wn{�;C��dkI��횞��]��$�i��
���>��I��S����'�q:��>����]�'|�E�Z#\q!��~�@+�TH{�7�FV���E�T��u6�*�a��ѩy�m���t����f�k)	���Oݡ���2;��(�L�=��}�(�v�yF;N�}��a��w�D�Ƀ];�DG#m��RK|�z��^�m�z�g�C���{
�"��t>YJ`PrJ��*�9�����m}tR��ڗ'&�j�Gb�Ag��?C��5פ/�!1���Lwp^8�`IT\�x٦f��cQ
ąg2����)ٰ��4^K�{�A˺p�,hB�z�!Ƨ����� �<��wf�"X�����ِ����[t��Ӵ	n�n-����=��q�|��bp�C��%�����\1��9f��@\��K[V��G��	s���&1�GC1+ST��z�:�XAZ�o��\�k�Ý3z5��N�f"'>�R��- 2�����m���O�BJ�$��3Lr��b���7�w_H�d���zҸQ��ՆQgQ`J��p�b��va��ºU���vW�J��XM{�4�P��*���y���x�'i�Nqh�T�:4?�/�������Q�(I�sH<��b����DH��K�����70P��Cc:�ufVG/Q;	h�^e�g���y-~�����"�I>^˓%V@|n��UN��u�Q�5 �<FhF���@���|_d�r{�˅���+K�lwNp�����_��m��B
؝�\8+�@�:�Ń��2�\+�&v������@�м	'A�%t�hƖ��S˷��zJ3���(<��A�~���6�umQ�aJ�Fe����<j�gG��U�H{�n]�b��rR�%nMޒ�;�X6-u��uE`}��m����7��Q&y��o�1Y�;��dT,3���}�ob�Gp/U�U�+P��ٿ�{ER\��Zu���Mi�q��φXt��w��� sE�bV�T �F�ц*��\�Cix�h��^T�'�g���C'o�~^��%8���B��_�$�lL��	�0�Q��$3����ө�P!���t�}�}?'��4s��H�sS���:�΄쟺�!7_@�2ނ�fL����XD��]���a�s���>���'�v�B_z����X�_�V��Д�֢ |\�\���!�`{Ώ�+�Zla��O8R��:3�/3��p5f���={{u�#=,��ūA.E����h�H.{�����g�ʵ�٩@�b���*��%o*8��D�X�Kd؅9�K�R��<��H�/�9hM�U0k@1Q�^�┱E ;cP�,��/���ٚ��C���/1��b���}���NL��$ǧ��){�Az�E�-�z�89�!<��(Z���K�0�1LA(�D#�q���T��`q�y�|����Vί�iH)��F����I���DN��Y�ŕR��h�3"����_�]4��N�`1�.zX��c�u��{1��\�y���ł�7kt���bHǋ
���Y�Z������.A�8���+|�'B�c��N*5����	;���2��+a7�c����(�l�y����QX���b���a���Xc5��gx ��Y?Ӫ[��䐱R�<4[�\�5>j�_R��@�sQ)��M���+���[8�eFz�5ZX&�q�D�?׳�.�y�qM��Q�5�ՊbvR.B�E� ֵБ-����gH�<�Q.,��ڀ�̭C-��J�O٠�&:��"W�5�a�@-ͥ{�o�|UY�頕��lk��$���+E�ۄ�=|Ț���0�}��~D��Ѽd�Ia��>������v�u��#%����3���=s?��O�ު;\X�*�ɱ�>����r�ճ�Hv�&&n��8t�f��C"��W���_����ZѫV(�z�q����\��0S}�/��-ى�AE���;Z�#B��_N<�S�4�ZL\T���WS[8M3�]��eU#�	v!��h���"H��v`��MU�|U�P8дok~r��������B�\�YJ��@�Ea��i[�l&u��S-O�,G
nA��z덷#��{�>����l���tv��}^Q�so�цo�R��L��.�Z���1�%(wK�#V��ſ��9�Phg<+��<������ai2A��u��i{(�n��ޚ{w��!x4����s����+ܮ{Z����Ş]�����n5Gz��_�]�]6C��W�I�F�0�g�����R�C�{!-�����-a�`�ҟ���f��;T��OsZJm�4"�;c��B|]|�T�!'�53*�{��`}X�Nx+����+�b2΍�㠴��L��S������(�ؖ@)9��I�Y?��L���F>5�a��A��ؼ�^��5��}��(j�
�Je,���p��"|�1:7+\�~i�Ө���{e�0gr����%P�h���g���w��3T�� �:h�J��NQ驽����ה���Č�֧�5�!Ib�R1v��o��q�gz��I�ݍD	��+ғ�@ˡ� ��1����&;�Z�r�ƛЅ6��U������_�^P��Z�^Xt��:�v!TRe�\%�gf���U9G��.��^*ڎS޶�V1{����,��\D Q�h���k��p��؂�V�a퉶�`�Ă^V���f�[�a�gσ�R�Wƚ��p��qR��}��y�^�K��e��IZ�k�I:/"��b�%�d�Z`��'9���y�qJ������������N��*��u!�9g��J�%e�>7f��&�8K��Ϧ��%/��(�E��k\��T��)��?#xڅK%��� V�Ov��Ӡ�c�Wy���X\`X�5�ДO�T�o.d�ČQX��3gqX��D�&E!C�أVv�r����=<����j�Iܽ��Megz�3JB�����O�#cA 	're��/�B��`1v�����7L�n�A{>R �yk��1<� ���-L�7:9�
K����6������8p��P������/u���_	7����b�im�٩�1f� �F3VYK�)NQy��b��5��\$^��'�e��%˸!J��C�G�)T����9�������d�m������!9�BS�P�Õ?5G�\w#d#HP�^��u�n��J�Չw��������мA��ÖO ����r����������`��Z��K(S���;��ۣXKmֽ =��8���pvp���^��wHd�x=sf��6�A�M�J�/4
�	���_Uj�S֔��h�Ǭ^aW��׷Ȓ���q���1�;�O��C���w)�@O`9��1Hi��|_�e���V�SfԱ������6X�5�ӆxhSN�Q�WH���?(��x������U�!�cA[����,��h�0��/.�~zV8������,&yv묢p�w��0�oM�)�\J�da����[��隦����@�H��g4|��	�3�����Y]Π����ym����b'��c#������7W�,�k�w.N�����;�H�tz�oܦح����>���s��DW�0�e�f���7�{)N7p�6� /l�R>W�0���%O�>
��޿�ͧ��1M��C��l�ᛒCb�(Mf`Q�Sl1~<�����)��ɹ���45��8 �QM]��B6�I�i��k��Գ��([S��м��l�K��A�1x7�eՙ/��<$\�e���z�pF3�q�=Ek6MR��7��>���ω��*�k�د{
t�8��9:Zi����)ȯL�,��`�Ut�i��DA��'[�`�d|iq��|�j�v!�=�N�yMNz�^%�j_��H��l�8�	y�����A31�+���h@	�{eQ��Q���ߥ�?]��A�M���7	����=�	��T!�.�ᬗ�!=��n�a{�����h�䥴QO�Y�[0H��W����0Ag�*>����eZh����p��[�;�n���C)�Ay#3�=ۍ���U�N:	��O�����qN۱�:���M8b��f�d���&�� �w� ��n�� �W�Ԉݠt��r-T�{��_��%c�W������6L�W��ؽ1FӋ	%;�NB(?b��a̡�.fUD�J&��x���-cm?B���"�a�B��՛yX�{�4P	i�>���ot���C���.(�N�k��E��N�X�_����H��P�2�c����+��" #�b����� .�ډ���En���#�a��h"�����6#�=���E��q=�Y�~�D��u��<2���>ݥS���hَhI>��{�6�#��yH�c��d�
�ӵ`BW-��t��
�@Ɣ��B����%c�T�C�=�g���}�Ժɹ32�.�OQ�p�c ݗsߎ�46͈�.���"�a;��m�'b+���Ճ���t}�7�
�RP�)g�j�W�)���4�g��ќ����D�����S���ǯ����A��YuN����n*Λg��� !��-�D�e9{$�o���F�HX��h&��^�w�p�I��ͲG ��{�c7��n������(=��nzfhnJ��A�Á�;�&���*I�����K�p/\`��ɡ�#�u�b< �/m6�&�D���eG�!/;S!gY?���Nt��B�o�2��*�
u3^"�9h���<�/t'3=
]��w�����)��E����ŏt�C�=a�L�vD+S���1��dd��H _w}Wz�pz����؊ ��vD@�H����@#��-C���4��/o���~��)K����3�T�L��� #k�a�!]a�L+��vaG� � t��۾�ʩTU��5������:�s�����,���pm=�St�*�����@�����f��F�䥉�cvv7��*	�R|s��Z���� �X�JۇZP,Ş�!1��)z���Q���OI�69�ڃƓ��ߍ��X�|������)ɀu�R����G�o�(�̴�u3�-�Jj�}�#�D�����8��jki������Fj)�r�"U(�tf�)���se����"���A��N����B+�bg� ���'Q��6�,&ak�q��=Hr��5�i��
��T3͔ |A�Í�8�κM��wȃ�D|�-A���
��L�5�
��LN����N��2o����SG�g��)^4����f`7���-o�O�]��9|h-��}c^Ôg���+:��3��� ��+d1l�ы�.�C����X��NhϾ����D�����7����w5�H���%���	�(�l�d�TIKQ�7,�;J����8ˆb���s��>pؚ��n��H*5��*�q��W�����l�FQoPx�k0@���u�	A2�q��6/�u#�sF�CӉ���k��nR�����`!>�,A��L�4�����7�5U����B�W��rw۫�$hAd��q�/L�Ƕ�4Ck�Fۻ!<�ޫ�O���k����8tK������4c���j*H��8��9��B�_�2f�A����^4�g[���%��NjL��F����j�F;�}�o
�?�Ce���I�T%>_6tk�do7;MήQ�� ��}Bq�L��]���]y�nz�k0ɪ焉Fmq�5�J����^����zQ0ȇ��C������
l ��]S��^����k齛���G6ȯ����,�:�I����-Ð�ᢰfxޱ����:���J�߲�����z�	�Jd��g◕��d����A�"�&+��'�P��-��Qy�-��X�x-)2��i_���/��B6���*��v�������s3A��Q �|�p���m�L��M"B����A�C��i:�����L�=���DH[t���@_��~�v6�rOb�6"R�N�ۊU��oq��M�	y��ӿh��>A������`x�=�u�"<J�`�P�{�}��p������Q#p�r�Z#���.x�z�}�E��L��:��)����� �;�������1�ᠻ�4Bz�Xˁs��X�R��IzR���S�x���_٭�W��U��k�D�2O�7 �)�j�t���v�HHR��⅑H���@g�C���*.ڻ�m<����<����X.Mx���Q%��N����<���{.`'��G�����Lgm����қ���g �)Q�4�_ެ�+���v��E�9NWlڻ��>�quz.���x�����x��d(���vs�d�9���!���Ya�r�T|�qϚ:�K-���-6=5s.�U�	-�Z�r�1��ƉdVπ���*��<� ��S�*��+�������불AF�-ԯ_m����[Zf с<�Z�ـ���óP�Xށ@�� ���mĮ�E��${��a��j�ce�Ղ��?vE���8���I%U=��<�ik�a�0{�e~pC�;V=	b���蕌�ï�~�k;�Vg��g��s�<]C{a�\˞�lc�W��Kl�@t��R+�%n�+}�����7�K?V���Sy�WDU�lƷj3r�h�au��=!��J[ ����
~��������b+V���E@�}��}#�Y\�P{�w�a�j����I&���DwF���~�����`	���YHɯ:���V��������D��m+2�ݘ+=�&@ٟ~�ߣ�Ӑkr�K�0��j؀:����`�m�k��ܜ1��hz��]�Yj���P�N��D��x~�d2Q�g��QG��-t.�Y�"W�-�gⷮ�-v�(���̑�Ψ�-�lj��䖍y�^�!Adю�4����7�t���3�W�	�xS�����J�bf�l�\xfzJ�8�.̈́�2,-��3����Q��V�`v��A%����gwp�ڻ��oe����:����0מ�b�Ӑ�/ �vKk$5���gQ���Mj��~]ì�/�SMqJ�>���9~ҭ���U�;�Tϓ�b��V#��}:��K@^�ha��N{ʋ���n�(a�l@P��ʹ2f�
@6��f�|b-(�_�b�%��qU�e�T<� rs�2�TO���x� �Ц�&ft�vzL���ժ�Q�_r_����X��+3�6��q��cy��(��ԁрU���/�2̆�ǋS�h5�@5���D��N.��*&�cU���-�U�`��{�V9&�mNVP�3��	9�uUIA�*[\dq����j��D���|��DMtp�-gQ������m���s�c�mQ@��uxa�qIN�&���+����ʾ`�mh��j#�B��V�*�ۋ�ԩ��������ǂlxO�&(��Lz�#s=p��.�n��h�_���EA��,�n�9cea߳#� p�̕���;�q�#l���*�) ���(.$EJq�����B��ת�㰡��y��8��T�s�.;^v�S�l�/J��6ز;�8ñ5傛��S�%�Mw6�3-�]Y�n�Q��BΒ4����- �\A�@
��|e���O5����t�:����%W2�m��^�Rث��6b�ec�y0J�C5���f.9���"N	L��cZ[ci���F��o����Ȯ�uz<O_��� ��E���g5BL)�Ed%�Z0�G3IO�*FD���.��R�s~ N��m~�͓�s�-�a�w1^�{�ض���15���­��kX����1�����GC+݋��t�7A���0(��s��:P亣Y]�'L��6
�O��U���cw#�̢A�9�=���H焪��1���Q����!�p,�|՜ 	_�r�'�Ž�=�$�����g�9�u��ٵ!���Wdr�͐��{r���W{z�ce*�q��ߗ�v$��+�����!�����C���,���G/_
5h��X��ʀ�ۨ��)oȷb$ ����0:�fp�_��iP�y��*�@�P;Dæ��_N�����>��c��v���e<wk	���N���E���p�{��G�["E�Ղ#^Ժ**a����(��R�3�7��a\�^L��s�N�m'q���������f\�A�z�����Cz/ϥ"D������c�.���\�e�����T�H����^��xSB�8²`+��w���,��<9=�k�1!���nR���Hߩ/c���DH��n���3�$^?� [,�Ő����k�Kz�E�6��5�����7��K 4���	&�xE�;���:��c�C��5��{hyT�}�sL�v�zʔ�Y��ߘ�����ۖX�G��}^�5�d�|�ov�qm)�bAe9�i�J���N$JE����dt@`-�C��f�r�?<xP8P�?�����'{C�P�z�i���ߋI���U��D�-�将v"�!�ͧ}͉�z����5$4��3M�|��
D+^�˼�T�S�S���o��^wOh�����G��^#-���l�ƥ)������Q�:&��vNz�e�	�s�-�68Uʐ=F���c�p��ay�0�NB����b��&r���^i���LI7S��$c�`XFzBް����\�q$�-_;vk@���^�y)�G#�z���+�G�	�L$���9�ɒq��߫D~���Q���H�V46����C�G��J	N������ �K��8��z3�	Ly�Up��r0�sNW:\� ���Ru{)
I�}�QۏdQ��.ގ���tvFt�F���i#�Nz�6���O��Jc�~L�=VK� �M� Ǐ��7"�T�kcw}[	����_y,��_-��F�j<����w)�Q���5!���:\�$%�&��3���fd|>�:�	l6_w��2���!��V���'S��y�~�tyV��g���?8٭�F#A�K$	���\;<��{��;�2u����LC3���H
Q��|o�tE��T�Sq�����|:�XT���*��U �Z��<tW��,�ŧK!����"�Hp>c�:dY���[E�%}��\Y*��]�'��L����j8��Z7qCo�!�I�U�O5/��Ո)cs��)���ݑ�t�cj�ɕ�k��?�!��z��G���&��u�!����6[������k���Fa���y��f��|��퍋�e�c>"z����	{[M��T>�  O������Zþ�r��F���p����p��OOA�F�sr���I]M��=d�e�$Ӓ�U[p����c_�r1��ӌ���IW�'���NPg�$��식D)7����D95lo���[s�$vV�zi��:de��7���PrF�?ը�D���Y2�C�_3���SD��3-�f���z�n2�9p��mMC���ms�$i�Zג��%�+��c �M���eYv<H�s�Ki�� ����)�D܈�|��;lmlR�>z�o���ԏ���m��Nm�TΛ��>��7�j���^�:~�BP6#�S�^�<�Lq
P�'n[�*"VW� �9���;'����.�P�Q����
�I���L��g���>pPs.n$AY~���{�\���Ɏ=&$�sZ��O#�s���\=�1�l������w����Zm�T��/�!�q4�-�#�R��[�� }O-2b{�֖��Gh�_ϒ��U�o�z�R�W<ԇc#Q����͵r{ڭuP�V��a��.�n��=�=�k�z/0����`�K0��ٚ`:���$��G��9W�>n5N�,�oC�"� ��~��&����fd�]�jWUȂ�==��w�2��4�@�t"`�f(��}��0�S���\VWpJYt}�~����/eG����)¯��hZ����9�B(5ĸ�y1�0�3��|`wm���ޓ�D��k��$��~B|�9S�ӡK`��NT��`5�K��;�5�m��>,/v	V�q�6r/n�϶H�,�:��Dɏ�������-}��R��}��))���P���]�����J�,�~cņ��`�aXV��/$RMɻa$+G��>�M�Z4��l���H��-���ζ�~<�d���jc�0�d���j]�3�U	���q��s-�.�C'�H��v�g/���O�]A��he8SRؠy<�4&s��Y���]*�H��h?�e �:�"�)9�#�uG*pa�۽D��[-	���I���0���L0�Tќ�9�%�~v"P��"����i�f�-���X��c�Ggt�6@�h^n���Y�1��'0�Vk�[Ӌi�E�"�r=�n���5�������#ү7�"�;���Ah����ɗl�Z�8�h�y�*�*G&X����M��;D���1����y���� ��N��t��D��da���ng���I
S�cbP�:	6�>;�( S�
�2���ݷ�s����%�v�2�^Ѷ���Rv��
�Jwq/�����QRr~K!����$���9��LH!�B�W2��q��F��iBf��m���9]��[�Pe ]�,��)�g�9��>�!%�d;��
�c�h�f�n_
�a��q�4:?���e���3|Ê�~�8CH��b�%5���m�����7�J��(����קZ�P!9FI�-�DR:��|t���_�;~˱s�Q�(	xD��[qD������O�P���Dpc��yQ����1P���������0znH���|A���T-���pG�@,��c�d�`�w�(u��!^��a��[�w�7E��8�.�����tT|�3@C�k��:���$T�r>R�'k�H�0I8��P@ y����[]�zQU��}>������w�bFy�B���
'%E��s3yKÊE�Ԉڻ5�&9y�*g�^G3HD�����?���&�s��.���^���&�������B�!�`裀q{ ��2��=H�x��f���P%V�!E��F��&��W|�7�ȬH1=�È[,\��:�k�NL�Yx]j&��&c��m��V�����B�Z�uBǢ=,�3�@zI��S_j�~[BMQ���&�$�(���#8z_L��z�p��&�!�1�-���`35T%��5���͒L����|E��ժ?U{�C�����;R�����z�U�kA�UW�ǨY �g[)P	�Kr	���c=/�ů�ne����]�SR�*p��
N�J_z/���,W��[��tѲ��^Ǥ�D���٦�=�j�6ύi4��t
=���`P&�d�̿P%ń�c]m��u7��b��8o���D���͜S#���19sy���dÛe�iP
��H�g�P?�h{�9~�l����f��5�xIF�u��p�&(��(��������� �g����/q���e� HC���}Cͳ �v-����gޭ�a9c�$��<����b��h;VE�Cۛ�2r&dJ��n�g�=�B��e������G�#�J�N�U�j�i�f�+18��p�Zi1��yJ�(�D��s͓��&&wwOs��Ȑ�Ϟ�q�63ᠰ�]�\��4��Ceo���M�4=�z|D�9�F ����xv֩�$���B�;�'���mԘR��	z���lr��3�y�u����M;����jaV��7�&�"���F�U�,!�7%����Ft�_o�ѳ�-�� Ҳ��X2�r���tS;wV���ݙ��-"XT�.�2�>a�}�	d	�S^��X�ň�}�43a�rۓ�i\c�^@�~�a��K���L�R�}�{tL+�pI�� �j�5-�GHF90Y�-����jr�K⫇��,�X3F�Gyd%�����U�����ʹ�p������s��d:��5�E��'�k״N�($S-�\i1y�h+M����l����֤�$vqz�Y��e��;��;\�u�FY��:�u���������<��|�M@o�옒$����z���^[ 2��.'�F�3Ń�'10�h^�]�Î2B�7�	��>�����,���*��0�l?�l�ߞ����2Ց>�ِXV�^Q��]�q^RZ�=��O@.r�[�c+�Bɐs�j��� �����] 
��}��K�l;�hCSD�b���D��|2�Z]F��!�H��AE�?�l�Ǧ���d�+	����"�]̲\�����kq�VH��F�z��q��E]��U,a'< e��Rg6�\Kjhy������];�k/2[�!Z�d!��n���xAP�f��;�"�=�J�t�h%i�Wx�PGtb��0"��jV��J�J��EYU�m��6̫i�����Bl�7G�٨ ���ώ�G1$7��Q7���i^��qqj���,
t�Ȼ:N^�UWҐD����N<�<݌�%�����"�_��F�<* ��u�\r�zp%p�U�B��ko�H��p��)m�!�$��I^ś��̗pW	�C��(#���c���ep�դ�ܮ�]gÿ�m�+':��^?TE��JĠ� ?�D�h`#�-_~�%�e��ߌ�"�4���S~��0r�}>�l�|�1)�:�Q�����5�����78��@��&���������F�GA4�7�E
�b e����?�J�(��ՉK��hܚ:�83���&�mo�?�@�H��1����C���1>AP�h�������Zl��V�ݼ���=�����Õ� e�K��#w��̼+�a瘕jX�PRVN�J]���[�w�E�x���u_�����Q�M�A_��\�;�ZL��H$�0��i��En�����]��`��M���!���8.`��H=�����Y�}�Эڌ��D�y!�{�>�1w��=LR�D#_�t@�1L���!��-�PS�P3�Ѳ�xo_��>,��^3������~�����N�RDq��e���\�w��W��hwx�����	-��/�,J���k8���h���<�,�a(�I%�F��r��x�!��Y�c2e��	�[�YY��}�hqXO+����:
�1*d!]���}9{'��}���� 5�F��G�c�7���W�nV@������[�&q4�[�R�L�#���(�S�Qf�R�K]3�y������bk�;��F8���/�RS��ƽCV��-_L�J�)�	��3
4R���<��µ��&hA�WV�.�s��5�p�m�e�����9�?�dCq���U�Tc�$�y=P@�"�AHGDO2v�ދ�Sn��Chx�!�R��-;!"T�	%H�z=�,N&�E�����p�;m�%�洃!���I9���Q���JSv����r�Ә��w����EQ�����"���!��J��{��V�}K�_�N��>��������5��]����B�y��i��0K.�m���ّ��PZ�o)É~[!XR=Yp�;��5��j"Z��2~j.�sl��5��N�e\Pl�ebHO+�����(t&@4��n��7��2��qQ��:b?�uK	��|�C���j/� ��"Dg����&�0�T{�%!�]7t���)��i����_�7`L�Q��^�������^Z�{Vf�.���r6f�d��B.g��&Ԃ��NT2{��"�q�yɢ�-e:�R�ߪ�4(�����ɔU��B7N��Dn-���Tk�&$�":�x�th=��љ��>�}	��V�u� �-�p.���%@86b��3� ����6e��<r���t7�晣��r�3�K�Z�CW��3xZi�-�9U�YDNH�+������I$��`���	�R�c�NDN�b��.x̿��i@�>Q����!�]���J��.�P�e���ES�{�L�)��X��V�2:d��r����H�6���j��ie�78w�N1�$8�����h�J�~Ґ01^�^AAi~n��b��ky�󪢪&����ݔ:�{����)�'����m'X6i����Y�Α��"�9��V=p�S������D�lĵ��G�A�b���m�뽣�m���VXf���/�r�4H�3�>�x�@k?o�뼖YzD!�ܴ)tt�������/�?�!Q\OG�Q?:����vц��
�h�I\��{�N�ܛ+Pl�+�E��e�ǋ��DNw�YYal������ ��wu!V4S��1�s�]s����v�T�O@��q��u}��z�N�!��ns���v$&� ��>�:���(4`�g����W��{({oV�bRf�"�oЭ��H������J��Gg�.�G{�����i-��8o
|�-�	{=�p V�@堞!Q:7]qD���TO���(������vi�M���cKG��� Zn��O�����ZkB�5�|���0[l�fK.�?�+�Y�h[�[���U�g1:��6K~���&�ZCL�@��BM_��u�h<��m�G�Ր�����gĽ|�?��f_�6Ktt�ڜZ)v[���膚YZT1����MKɨ�m��&s�e"�f�?(eD�겠����/,Z���[�Ϋz6���w�7M@5z��I�� bh����.��Oo�hB��;�A��.'j�Tڟ6����]��h�d?��e�țNw(|�Kfm[R;��K���Z��D����ٷ%}��Z�M�QG���*mW6�:�CH�ՌFZ�Bk�;ȇ��
,�Y1=��GThf�V$���*o�j#�T�8,�)iƇH~s��H+|"�>��,��cD��"�j�}��#&�\#}� �� ��P�U�R���t�j�cڽ��D&3&v(�A�Χ�XJ��T��0T0�\L�v���/��M����m'Q��Gy�.�j��"hb�4�t�� �����Ƹ��}0�h������hw͹��!5��#E�L�D)f����'C�	�v��	�i4l1_�hJ��x	��o1��v���F�Em�5td���qt#��a�[e�F)�}�j���A�d��
�s��VӺ!8q�Dg)p��n��(@������g`�	��It��XNYʋ�3���չ���D�bj�'�	�Iy���#1�Q���>A6�%	,�sg�� W]���eP��j.�:%��r\�NlF6�-�iN������rZ��F-&��������s[Y���4w���8~�8:�K�l%��6��ꍌ�ӍSI�A,���ꮟ�e��$��Z���L�V��� u����'.jR�EsչC=�����Xj@����L4J�#�jxZ�+�Ef銰_��z���ɖߝ�8)�d̍$��?��.&���5T�5 ��Jo��2��o���r h�a�-���@�P	�M���~r�6�T���,V�s��^q����I=�7���D�H&˦̢(�B����o�D��5��x�zQ��dQAҚCu���ti��k��T�"*��r��"�M��!�읈b�
�Jm�F��nB&�C51���~��/�)�n�������6��L�$��ۘ�q�`�3=~ܬ<o�{�m�j2�J�;x�?�,�α.��5/�'��YUZ]�����6��-�u��O62�K[^�:GWPѹ!t�l��������Z�z=_��*��ƨU0���]��f��ꌾ�!�ʀ,�ҷ{�`�e.gGQ;���H#x]D姭Į�atޖ�����Ϛy��b�70=@��+J�(t*߬8H^����$>[ΨT��Y���$��	?.Qً<��,��+ZBU�ڴr���˝��K�'���اC���r�`�Ҵ��1$VQ%�Z���������<~�#�=����"2��y�4h�� B�z�"�Z�K�#��|dj|����[MV�7-*�_J�����C�>�ZЊf\U~bO:�N��'?��ԐL:���m��G>�U+is�SÐ\�қgs�}�p?��������9��$������y��ↄ��{j>H|q�#��y�&,	��<��_Z����~�F���F�g-5�� �XW ~�2-_��݅����Β������JXͫ�պ�>����#g�]ζu�+ֈ����[�E&&�Σ�s�hT5J�x��AfK�%�C���撕tDx����/L\!�$������؄����>��tXD�cvGV����S�*���V��`���n�O�`d��,�q,�	�i8�$�#�|��:B�D��	��D������D�j����N�3�r�_��<ge��Έ¾|E�0��Q��ns�ˢk�u
�����Xl�ѯ8ZE�U'ʎ�m� ���,����t���N?3�;�I[MgD0�ِ�4!�>eg��#��_E9�a��3H���A��Դ��|x�onb��:�y��ۿCJ<+}��H��io��+��+�Tx搩���r�<��+�O�5��9�ǰ�I쾱d�Քa������)��76Y�}|��SŤ�r!/���v"��3
��f��?�F@(�|����kE5�/d�	g4��*1��0m\�[4C���͏���4����$F��MdF�x��(!	��`FL��aK!�o� ;U�=��QT�ԁ�%��*$V�yqD�~�$庎X�"L�S�ܠ� ��&��X.��!YϺ��|�����v|�-��Tco��񠅯�g�?{󸗈��588��v�FQHI�#ϵv�#' ��<���3R���2�)�M�C�%V)d�����zM�u�Y�Ǳ�����Y���5N�}&6#�7c|�pJ��"44�jԂħ#-�ôw�1��c�g&E,8&�i����M���Z���'g"WLp}ۧ��ܽ���T���SƄ�?3�����jF�xiB>v��$�Yi-�g?OhyZ�����n1�e��mC�6�ZW�$N��pu����)�j�ɨ �x����b��}y_W�w5|黐R����"��=:��"%�r-I
 g��PG��	��c&W�m.�Q
0���|*�s��\2b�� �$�L$��#��/ԙ���g����4"[A��?��*�� ���k�����S�Y:�z���@:��һ̷@kv��0)�Z	Aa��+�o�9�{^�!������K���|q�7`�G�[�(�Mȏ����.U��թ�ҵRIE��A���T��L���y�+M���=�ƛ.ϳ�G�~�^
C����R�&�S9�0f��#[�^wt�B&4���~$��a��mf���_��Ø���D�`+��������׻�<�1<w�X7P��^}��Xw����Kj�&�s~fyS�١��2�6dE��^$ߙM1� O�O#z$3>��WQ��;��\P⦖��޿Ӄ˿?�����'ldT��B'Nm�N��p���� ��`�.4,�2Dx�����:�3$1�$
�c��k��?�v�@ɗ7Y.QU��IY��])!�~�Σ�#�H$�bp6y���ʘJ�8��u\B�ޞ��m���	�A�}�2oq���1֝�O�q�c�7��� g���s����Y�����@驯H��Y��v'�q��-�D�OP�Ѓwt(�<�\A��?��61�����L�e#,\'�����F��K��$G���4\�/$�f�t3!�oR����J�I�x�.�k� ��{ń啁f8u�B*�9U$h$\��mGn�i�v���8��V�F�ܤ{���L&p|+?�)��	� ̓���,4.�@~S�ײ��k���Yu���7Aap�vn�Mx}z�vVP��k�BΙ��4��9hq>�פ�I1bP;^k�I��OKDT[��E+�&�`\U+'v%�Ќ�b�6�]�o�T�Aa����*i���O���6���	5u����T\�T��%�0�����l�)�<�2���Jd��������S�{���W��[�9+��2Y#C�k�.d����ʗo�����թ%��!�N�8mgT��(*���š��$w`���
.GQ��C}��]<��}��'�%Ҟ��1���)�4�����i�Gm�u���\�'f��j�����^SR�a �\F�����0v'�]~���(����%pR S��I繣�Oc9�{������؃j\0.�V�
}�'g�І�����4(<��&!�p��������F�aV�W��p��PӪ1JD4�p�|A�+}0m*ѷ�'t��~£կ��t)[����_��\�_ܷ=���%H��a}H��^����	V����o����G������x�.�]�ؓR�7,X~�.�D�?�v��ll���OK	�*'���d�JbHX�OE��!(��>
bl� [nw�Hwݤ��稂\L�8���6>��H��i��U1�$*�!�k(�d#�1�͙e��i_�æ��o��D2R0����zg��2˨Kˋ* ���˛ā�����W�\�V��:���]#�Q�N�Z3��������O�Dr؋=nR�X�Wb{�R�Sk����>A(uW��eMɦ+�.�-�, �;����-�'�.zT�3?H̰�)'�U!שp����2����bx#`���.B��%�}��T��C�,�R��41t`�s��xÚ���|�ਁ���n2��k�(w�?�Bߎj�FJ�-�C�aN"n�#(�%l�.�	����?��:��yw׃��A��UH�uM*J�/Wj�H[�S?"����([;��9�����c$�2p�|Mo����{��{;[�����h�����ڸ�Z:�m�,��k����^/��<NBEfZ�>���(h�A�;G����۰}���=�s�o爖��e,db��?�I���2	��-�"tJޠ��@g�6���ҒkG��V��i�=�t�	ᐧ&�g+�ԶZ��x��D-�en�zf�`1�C/�ô=��u�"][e�q �k����5�������v�hqr��^ٳx�U��|(d`vێwԣD*6)���#4�IH�W�,�$�Vm����aE����uE�q:iο�N�Q3��Mm؉��ǵl��սj�*���G�>bG�-�͠�d:�Q�u��y^��v��������o8�wlݜ��
K�G�HnM%H�(�9c���9�3>�(T�<���I�ч{���9���c"��J`u��g�h�1K0���)v��(4�I���mQ�Қ=��PY��31M����pL����a�C�C���x�Z�F��(���&�]�35(b��mU2� 0!����nw�h���M��Y�j6�8��Xf���Q4[t��6����Y����_!�4����^,���l��l����LN�� `8��c�S�)-̛Z��ϣ5��p&|U�!�A��Yյ���x.M�f!TF;x��+�e�e|�ڀy�M�^����r����+��[��P`�;���S��
��T��4�#zZ�����%���|����?D��R�61��`a�.H��@:b¸��#�㭂%�v��]�u,_���hG&Vaa�����,�6j�}u��U�9�ڊ�:�!��āg[��� ���JtΥ�I3+�*"jA��P��/��Ld��);�0�c���w:B�!p����N�,�]�u��G��3�rK��-׉bH;QMu��e��1��/3�͇r�������'��<p vГ��_�AAJ#Y�%a���du|L=��U�/p�A�y�p���H�Z�U%?j��Ä��������pS�/�^�vJ�f5G��F�b�|b��,�W���+&��}B��M���HA[�@��|;���Glׯ�P\p�nѕ��C�������hM3���t��k1%���we ��IH����ݘ�C��r-��sr4FqE���;9A�DlhK���t\�$���OU�l��{pgQ�RR��	�ҹ�7dGu�3�,&I��#���Y��ƈg"ULqFnu�&M}%+m��-^`�\�1y�	h����sln�*6���H�]&�G4�+h>���C}��n#��漙�����ƀ�$m`j�8���"�<b�`�+_ӷ�W2�4��{U�m;}ϛBǄ�j�9��'����j��*��ɵ0�A�zi��c��y0k��}w���>� (�`�r����c�K�A#Sگİ�w�1���ϛW�F������]vyP�⧔䰇���D'ұ�Y�	IZ��$[�k0�SXC�!lu��X��n2�Lw�.w"�G�̝4&�5Ay���蒺s��s�- p*��{*��5ڭ۸/�n>�-(��K`A&%�����,K�����������
���3�6䗔�E2�F��h�͸6���|�l���'����OI�hb_u5r�tC�ef�:�z��� .M+�R�n�k��"f��T,ǀ���f��;#����m��T'�z0��7�ǫZ&5�C	�oc��cD�T�	Z(�^A}���u`L��̋���Da���je�@��d�j Д5�@h�y�=]S0%�?�h�!-R<�{	�++n��?���KF�nW�ԫ�wmO-�I5��%�����M������2���D��M$���{�^���)��U�T_�ү� 2M�+wx}D�i�D�ӥ���'i �W��2P[�P�7h�}u�S,��hO��6�,�Ʃ�[�0<�m�@ɋK�!<�С�^�k��:�15����,����������؊�����vۀ����ӕ�_��r���z������|�R&+:�$���Lh�sG�L��0��>���ܐ�#��Ή-=�w,���U%�
�T��iXި��M�F �%0=\ؐ	�O�hq��QR��CFnʙ�4�0���*��qX|�:Π(>n8���6�)�=$���j�	<}��4�zI!5�up�F*��I��c�����3L=D�x^�+]�s	�}�t����:DX�N��:������a�t�1
@
���wA���qW� ���<�7��e��7s�K�K7 x��e��3O�D߅^ $D�ݿ�guFg[��gcxZA`$&,j�h�~^V�=�|�Qַ�|{�4��R@_���Ҟ��W~�1��_l�5qB#�*U� =��b��>�[;����x��,ǤK�����y;i�g������)�$fRiΓ:e�U�b�6{7�o�{1�I�N�%��#��x����w �(-����f8�2>�	��C���������� �8�� ���`�@aZI�u��7��E-�OŠN�gx�2爤9S��d�$A��g�u)ܪmS�0�'�	1���L�o���ݗ�����/�����jAfHd�_�=�H��[pO�N%�e��k	/�+U�{	%C=~�ݰ���Ia�J�^>#�6 ��H�o���CB�+G��vb��H���箾��7j�$�Ç#M�kL�)jo�Av��R���k7��0w��	���sL��| H7�w�K^\�$K>���۴��������NM�b�,����XjNS�;�oȊ���\�Iο$+c\�I��������7Y����9@rv|�ؠu��
ƃYN��΋��.�L^�]��^�@��	D/�������ރ+�x7c��6H�+��@��G�MAzWx_B/)�c=z׋�cy�T������6f�1���t"Rؾ9�Қ���RkV�V�R�=��Ҩ�cJԩ��a��S�q���	��-��N\��m�F��& �Vܠ�,^.�D 0��Q%bD�v/5֚���v����5�_�(�FPd��Toٺ�m�g���������S&��,V�9�𹨖� ܳ2�e̅sҧ�KD�64Cc�d$t �v<�ٹ	�-�Ī�؇m���E��n�v_���6����a??
����P>�e��b�t���Q@�peo�r�r�U�R	�-�|i+��|��<�cͯ��6�;�{m5p��~���oD�ʨ��_!������N�$,%��S�c�	�V�Z?�yD����w[�����㣼դbp�B�����~G�t5٧w�抑���~�+5iHq넭�����΢*�I� �)�"�}�}&�� ���3��n�g1 �.1� ���=_�������KXc�#x��2&�k/R��}��茸�3�#ÛL��g.���F9�IN9��W|��	*�Đ�"f��`�ޓ�ӈ,sG��I��"�6ռ'��1�L����g�q.}o����`#?��
咁H�AI{_Pl$�u'lKR<���(�{a�HB�+m�H��%���?�k�APݦ�R�� *�w\��/ل_w���]��ەs�]�g�H=��R���N%�����Z3�E��
*c:��W<�8�����N-z~Q��e�Lc��(1gݮE[�O�%v���S
���N�	�kmb���n��>+ܙ�J�q����xC�3�yU>����4U�#y�R^q w���7D���lq~�r��e�>�H��֏�P���P�$]�.�H�4�;剹�.e|	@�!G�zN��n���J\�T���o�Jq�Q������M(�+6%Dp�{�rs~�aҼ�������܍���E}�խ_�ē��p�ÃqS�|]F�r'�8�������jO�����S����C����++�� X�pbQ��$�0`�v���!=φ7I�/Ɓ��,�o�OE�>-�F�!�C���b�N�<��FJ�Z~���hC��f��j
���E�����|c �Ts�\�E���W����~��@�F��3�&���{
_Z�M*�.MpQ��yc��O��⁣v�˙�(��X�),����WM�ٱ%���(��'������X�ߚ�ߧ��}D�6������S%��Y�:;�Ѭ��G1�N�'�P���  ���V���w�LEAbX�~�dج	XU��9]~�Bxmi���s���-��"�����X���$�K��ya]wI�R_+�𙷡'���W�:�v��48���\�뛮W�!�G�Qz_�ő����2 ��ݭ~���q �O[�o���Tb�6q�
������\8V1v���,d����n���/bH�i�|�kn��+f�wë�j%���M���B'�20�tT��{Ir� ��K���C��i�a�Q�P��a<]���J;��*��oj.�d��I@��ʶ^`���[r�MPC}p�S�g_�	@�\��r��<@���{ۗq蕷� ۜY������)����6!p^d��z��&D�-������N�,փj�-�@խ����ºS��^.l�s�AU��	k ��קJo\!�v�۸�S*l�����@}�aP�ߎ���Lq��� 7�l�~%��=-݅�"U��e
E��&=}�uX!c~<5y1���)�eF��L�3��ȼ��j���k�^8�]WYW��S,�����]���m��.��^����?�K�#b����V���29��8��x۪���[?CQ���
.
�zY���)NnK����IT�l�� ;��Ӑ��u�����:�$Q�S��;%���n�_�В'��;�)B�@K�<9m����}%#n�3},����
�aRD��d��~� ���ĠK#:�v���T*����0dܐ�Sl;�N��E2���J}�Y� $�'D�h������]�;Fl��Hg��\H�䥒o܅M}�;Re�q���1�c}>��[�#���J��^hL����g�Aq��F^�y#j}̍��ߐu����Ke͌�D<ZY�ɴ,2(��e�����=��X�?v�]�Q��$zn)� ��Z[|YM�LFb�?�ra�!������y9>UF���W�HN6D[�hu�f+��a��iz�J|V	>�BP�3����H����ZKd���I���1��7u	�řs[���S"���z	3�5J��1=�(nނ2w�ɂ�Šv�3��]�g�G�o����y#R}ٵ'�?�u#c�G2r��9����<�(�
\� m�(�r$� n���M�	���-������hBU�F�D���������2����L�S���B������)��L�Ӿ��i�E�M�\� z룶V�B_f�=�ޝ�u�XKs�GA��؍um�ё�ԌU�E����?O�"��I�GlJ�V�e��v*z�X3!󜕞k��\�<�����͓R�K�+��ȹ�l��!���s�B!l�R[�����\�*�����;b���UG �ã�xQߋ�D��M�y4B7 ġH:�{��&I֞���k��g��G��d�P��
�MW=�j$��DY"f�?o�Bǽ�,��U��r��d4�g�A�m#��q��>븀+������l����)��Ԟ?�4(��puH�j�i��id+$�a^N}��V}k��鷖������U��ؓn>$�?m�1Jd�G�Zڝeאue�%�j��R;!���b�s�� �	K��.�(J�N$�э$D����~�nA���!�_U�w��"����1��B�bM���� �1)�*Om\:�Lb�E��&��$���x�@ }� '�y�U|�$<*!�����Q�L����,k�<�$[H�}%����!��K��ח���A��n=]Q�3GP����b�@�h:X9��0vɼ=�f.�<m?�q��8�jj~�XT�Ks�|�@v��j�b�5��Y�b?рI��v��K��]!��n���h�jt�w�c���]%�itM� ���Ui����wW�J�;��cՏ��wK�6Z�$�\"�7���^[�1���<�@@�9c�q�.�����"p�#j��9
⸕*C�]���������c����4l��Xc�<Sˣ.�%�"r.��c������͹uһ&��V�t@
	�0�l���aX��/fL5y<�[����'-� �� ���B$S��5�k������@�68��r�� ��>�ak�";8Uݳ{v"���Q�x.۞*�S��1��[���b���݃�������]<;d�F+R'V��\vЅ?��1#���09d�8��,oA �q���8�WJ�<l���s�8X<�_��{�ƣv�F���3M�/�}�i��c�5�w��OCC�aRZl�h)����ш��w*4f}��!e��&��	�[�M�?��+��:,/7@���4>6���5��'R"Ü����	i8�ԕ��X��ZF2((�f�8�V/���� ]�ۘ��|)>�s8@�[?{b��̔��W��[�ϝDE����#��vё6:�Q�t�E���`N����5�j�n>t�/<.�7l�v�s��p6�g�0�7f�e��r���ւ&k��Ɏ��v`s�RH9ή���j��07~�R.�?�D<b[s����G&�Ҡ�02�O�����cW�n��ա�2��@���O��3~~P�n`u�w!�\�{���)e�a"�d٭_Η�x���Y��^6���0��b�����ܗ� <�M7�h��(�zx���wjd�|����ɍ�'�;DE��B��� Ї�0Ɠ?WMKD�L��v���p/��ͽ�}���-;M��������tnm�,���O+
�/�<`nLu�tb��7�����C�)n�>W9�V��btm��,�ͦPN(�)��;�dd3���|�~����!�z�54#p��������G�Rz��ȟ��Ǯ΢#���t���a:*���F-g�G4ڗ�%5b K��{ w��{�[y��>/TKT��+ς�V�7�@.O܊7��^��eZ��'�Z//Ǎ���-��O��o9�v܎�]@��ג���&��|/���]hE������˕���ù}��ū�ox�o���a������kr�K��<����*�8�W6��Q�
����:ᖀ��fN��9��e�ap��]�R���ڶ����[����#����U�@��*c�>[Ew�O.�com{B�&��=u2�)�
T�hbs���<d?�X�x2,����	ք��d;��[�M��kˆ���W<%�u�.�u�ҭ��B���((G�ʟ��5����᭰�A�OvWC��[�I��`]�/Z�o���b�z����0$o��R��ښ�;��d� �n�ZhĄ��z�]�������v���V��mg��1Ť���x�+>;�'=�b�%s,OBs� �iɦB�v�MD+����y&�����pvvN7B�h9a�H�շ{7R~��^O(��,���G�[��*.�[\6����zE]y8����O5�H���mZ3a�� 4�ƝW��)�X􍢈��k���z?�a|�@|��U�����Za|Ll�,J����F��Ʒ'�g��%X��N�^c87=I��VA�2m[�bĂ����Z1�ȕJ=��ι�K��d]��ΌZ��l��hpJ���a�d�F�5�f�ۻͮ{� ��[��ԓ5�����K���x9�ɚ��K���Xq��W�,�G�O6�|�u�J	�s�P��=#ߪ���[��^�����NH���K;vE#q1
��Lj�x�6����Z�(�*����{��%R�*������!ڟ~�:�d�t�z���@��c(��}�@��~�T,��Y�u���*���g��~_��a�Y3�1y9���S��'f�`��*0�Eycc툍�	�E���|d���A���u���{zU/�R��/��5�ʕ�"�q�:ʌ�R�u�H*h��x�������3'�3WpD�4j�Ak�A��"�ax���zՐ0���/���|G�1}�;�_��VGu�r���������,w����6�w�k���F ��&B8#P��?j�Q��W��(���YĬ����k�0͑�"w�s����A��<��?�j���RCO&+"����p��<�ϘB}~$�̞���N��W&D�k�Z��yl@�K�����J�DL2��@6s��S(�c
i�?)s?���(�a��'�	&)��>b��X9����~-!&�^��V���x���y�^c5;oyE���Z�:>�����$M�q�t���,Jݤ����#�p��+w�w������I�Ut�9T�-`M3a�Q���m��R%{ ���F�l�Y��ĴR��w��ݢ�����P���̮��4͞��v���,�򘡴�Ci_����u�gl ��Z�b$`v�a��&Pͧhk��5	7����NC�G��m
�{	�����L�/X�6�x��0����#�ˊ:!w�]�/+�|��=�u9?�X^���𣋓bm�F�ޕZ���3T��q�~�-�5�1�i*
��r��MJ�;�'8kvsA̒+��c<B(LB��~jW_���
o	f�Z	�	�_�]���ȄvX�^���s���t]��i'�ޫ?�E�b��R'�����Lz*"��)�e����Re��וE`8U�b��b+'/Q�I�G�)��c�t;��/1��Wc���M��p}7I��"��3�1L�!�j�kA2MP�DO�0����s����s���<��g��������Bc%��F���6]�RR���M�����ѩ@R	ŧ������;������lǫ�J��^T�'�Ĵ����Q�s�:-}��Jg%b,S-�1���.�c�8W-��������O��"�%��"��f�0���ׯ'�Y�!�nX����� ��F궭Ͽ� ѯfZkBA��]�R��<~������ѹ,�#���r��d�����1aʂGK��t�6��4�U����~�������*/�ԋg�nZ�W���n����4�Jo�����г��X����Ҥ}^(�,)י5�tKrD�ڟ	-f=]֖y~��]H�`�X���_M��ˢ�,�q��zb@�ɒa���<�佌H��f�?qRgr�颴=���o#M71�1�7��Q�m�%M69:Ҍ�}��*�Q����LP\F �`X��=��KO�|!R�Z���%���b�[��D����խ9����y`�a��&�Ń���}׽��R�"2p��J��$7��8 H���C��%�E���O8����_��"�A����!�%���1
���o�I�Wq��;�u2g���<��8:{8�B<��w�f�)���L�����q/F��L���������+��]�}Pɻ|2��7[aSp �u�>D>pp�g�9�M�6�eJ��X��NYd(���p��؎xK�;��I�&��w؆�Q����������l���ؘ:J*ϴ0xk�Y����!}�تC�4�`��$	��D�S|��M�+h���1�@�ǂ;6&�Bw�����N���>��(��
�G�5�U5�H[���K��p�M�8,���[&�o_L����Om��>kn�Z�p�;�G'nS{�E'�Tq�ɤPw�N,E���m@p
e�k�)+�����P�i��:�h����y7�a[6@Ŷ��uv��O��B��\1o�����0�,3��x�*̰����)���W�Z��΅܀E��^�B��������(�=��4�ŀd֙��b�e�B)ϛ���s��xjRi�\�;K�im���=��W�yai��#��}�\	";A�uՇ|��Dr�O���֤�y��s�[��蕤����:��(��"�l�J���tmj!��n��<�$����u�=�]�*]N0�5��p)�˩?��Dx���u���A6ͪ����Y�]eָ� )�mޔ2@V�xԶ`{J����ˢ�B�����s<�O�[���l�t�}_-���s��H=� 0 ��� ���?W�����3��g\�b<A�v6��8����g>ϝ��4��[5�m=݊a:f��gT?��v��\���l�����fI�)u����#\Ig����W����P�>�5���a��_�%d3��^Gn�*#������>q�4s=���o@��2M-}����'�[�����C�Ui�����`];�x����m;I�ʷ����Z�f��[TG�x���|t�o� ����f�9���d�-��~��S �g�Y�X�1G}"�XǇ d*3�W�c������pq�9�7�~������q|�Wʚܗ鬓4*�B��d��wA �¾~~Z��CaD�P>=�>��DI	URv��9n�
L��ÄNN��6H�����}�SuK��,�x\<��K7޴�'�i <E��lP�ܔ��!JN��	��J��S�=c��sX���0%a'Xwiա��T���rƦ<Go���M��@�
::z���P�J���UE"����c��kI�y��_���n���6�W���w�p�Y3�('��v�w1>�ϑ��8�1W�>���v@F�Zd�"��ZUF�3�~0�p��ѹ֭���2Z�Luf��$*r]@�{"i�j�q�y��>o.�`��Ѳ8���������~�:`S��z�+�:��O��O��Ax�ʇ9S�� ���J?��g(�͓��$����m�K�#��f@�7գ(E���P+�$)�C~"gS �1�ϛ��.#��8�C��:�Mı���cM��2	���!˒�b�>�M���pG����'M�ܧ��,}�+�D���F�'�yv��f�P�^��E��u�ށ��(��z}��z?4}+.�y�6I&R�Ƽ[n*���;�L�};_����RѬ���h10�x;�B�%�y`Rd���=�����8z���{g�l��C76�����)E�� CpE��\��#Uw��yl�<�̍��cvl�i|]�V��(��ښ�IfC��P�|�?��R���G�oi�3H�. �K>��-=w����]�9��̼і�"���ШhM����g���\1kc0�ؗλg�W����joU��̶	�l	{F=)y�ҝ(~|�bb�F�ڻ.�
�������y���B# d�J(�ث9}��h������`�c���|�1Q����J�j��FwiK\��Q�r(Yf�C�3��c=��CB���2um"k$IE�,���
d,#'c~-j�[��xߚG(�0�G���%>L�N
�cHZ�G��h�?.���׭����/�}���RSS>�T� �Ё&J�{8x���3F��ְ�~��Cv|��um0��`n�uܑ/� ����?��O�	K���]�E�M�g7�^��v��	[@N�·��O�細P�4ử�.��U$VG�\��.%�f'�L�\ƜrxoU^G�L^�#��ZrbɃ��OeH_�:�L6�@0���o��T&yͥxᯔ�&2Mdg���S,sWE
�2��d!�SV�����t�>�9�ep�eC*�ޒ��L�@p|�Ӿ��1	7�z:%���h��䖍�H݋��t���������%9>��\P",�7��ND�*m�Z&��j�k��D�?���vD��t����C�������ص-�å�!)�q?9��s��̛pp�ض���S�c��&2D|�+s��v����u o��0�nF$��Y��2�a���`m���������>��S�������`D���5��%0�+"�|����D��D����G�x�d]�3~����UG풞$��L]��V���3��93F�}S�Y`��=�x��B�	�B�	��4��V���vG~��:���k��'�	Hp�Z�Y[���ușsR�3B0_���q[�-�@L��?�p�=W���\p��b��t�E6?����u%���g��!��]�d�������ڷ WjS\�[*�C��,4���c)%����Y`�f�TxG#�w�WWTaFF��G���Us��$�W��`�.!�*�1�T �?��Fli��5Pyu��p��uk��3��t�N^��
�PҠ���yN���k��'@3_<(��F3��;�3+6d'6�([�0;�y<������oX�%7�9F��9��-5��F��r/?Β�,.�ڨdH�E��<CD�&��:Z��i$����J{#�Q �����Q�-&� �&��}!�Ngq�Z��?��В�� &[0֙<�"��oa�܅@I�Ȇ���U~$8an�X�o�%S��aŃXarFIM�w��K®��S�D�{uS�@'��"ὃT+�!�tZ�ǧ��.8�pfU�4����	��%�GA�n�pXwh�H�~�ߘb5~� �>�:�!���6�jù�}h��Ak_S�����~'$�pu�.\���0������uB����@U���{��<=�(gՏ��W�+����ш���W�F��qBZ7);t2�ZX#ŉG�G��c�'��w`����Z�61F:x�@.����R� 
7C[���M��mj�P�u 
1��JB�'��z��"\��9�'����n+פޏ���p�di�R�9� �H�{ұH��pg���psqH��7����ɟb�*�1�<�s%-"��N��;M�в��Y��P�b���m�u=���/���qI� ��O����?���.�v�k'�拫E^3ꉘ��6�ʍ���h��F���2f�"8�w�d����T|�<�{u���B���C��t4�_(��˯Agz>M��-B5�!��vƐ1P6�,��e!O�Ͳ�H��r?b�S_�r\I��@H]q�.K�aX�c�!D]��u ��]��zF`�4��Im�w<����l�m�wUX{e�f���t0�B0����j�T���6 �W\(����Y:ƻ'�����ۆ���W�dH(��ϗjՇQ����l�'A��U*�Fe]��a���7�|ܮ8��[[(�@m$&�� =Hd.|ad����<��kQ�t������F�|�]����Q� y�/�,7|���k��+?��z��;�E�;�UGS͓�0��Z�GkD�D~z��=��ѓ k)�at�e�"&�Ȁ��-�[�un�Cx��ʪ�S������(��6��]�/Wqq35i��^�$��1}�Q��R��'������I���Od�>҃=��F5�c� �+�m��5��*ѭ�t��Ɯ1��Ňږ�������C8����?�I���3�&������N�쀣@o�l���s��qp�؄�߀�-�C|�y�8�8a?�^��=��.�C*�7��]|~K�ԧ���;��qw�j/���P��~�u4
c���K����S���Z��[��e��b��S�I���h���5!��V��� �4ǅ2wƶ��6��h'�|�V�	eQ1h�}��*!z�����Us�R:����GiϠ�$Lr�:&�F�����?�Y%��$�?�� �p4�s�sҵ�>�;%J@p]�1��N�øy$w����a
�SjS��[�a����^�3�ZR��K[7!=*i�_=,��ēZ�}��7���H�c�"���>[j�\�^����$8����}Մ����z��:���$����⹚�]�9�A��U���V#�G�	ҴRѴ�dHSӆ�>DW�/pҋ��!؇��TP�c+^&�D�|�>
�<I a�I�R�u�As`��t�.!�*�2%&�j�c]�i\��#+7P
�r���.�G�0�Ğ�땛�F?��%��J]���`��\��s+�ўHkh�M�E°[��^��P�C��<c��+��Lb+�sc���y�͜��tX�� �^�g|1��5�υ��N��AH�R�)���տ$6�@:��	���Ya8}�!x�P�.��&�<^��Y��5�E��k���-۽2J�����}+�k�N׺-3�(0D6n��R�z�IHq���B�TG[(��t��ݴ��\h�jm|$q�!ݻ7;�T�'�u,󝉵#�B��r�-���@b�X��7L��P��
���{��.:�0бh�ծ�U���i�7;�O�ئ�+�& H%��!��]�\�o9	
����N��9�&��S��8Qd�+�m���2���<�z`�uU�u�͢P�q5�������&[vn��s��]�^�VLe��J� S
���wj������TGxgfUG�񎕙MԊ�h/��ֻ'?�?�	`w�D�n���n��>0.�o�`�M}����]�8��5;�#�bru�1ÞʧB�m���*x�!���e���d�3ϑf@Z������#4�m�_M���!��z�lʞ�k6*-�����X+͎�A��-n6hsr�<s��!/�VI��D�(=A%ZMaۀVU����J5�n����9d���>X���!v�_%U����۫���=��QB�o�@�^~V$*���pL���r�2�!GC��RڰC�P}3�J����*�WTa;q��Ej�]Dx7��w��r 1�Eķ1�i�����'��4��߉A�$��~P�o��Q?��Lg�骫Ý�i������n5Y���{��mK�K��M(�A$�V�hca�����ߪ9:��m�We��t�)��Jظ<oj�<���X�%�9<���?,h����3��%����:K���V���Ǫ��:a Gգ|rru�Ɲ�-�����d��[j�0�'QL��G����BMy��/��z�.�LV����{�\�e�!c���e�'F�,�H1��^ϋ֒�p^D��<&�knm�o;�����B�_'�zq��R!����0 F������%�M\\���d�W��ka�Q%(ȚP(4���j=�&c��A����[�8��4�Թc��M��f�]�Qu)u����O�
z�hf��D��L���̮�l���$O���՘�i���6k��X8"�|Q�\��҅�S2��5�z�b�;Q�	"�R6M�+%&V�d<����Ο�4��*�!�iL..���jE �$<z&����۴=vn{�6�#�eP��	jU��/�Md�,��KmZ���8���;1�싿Իʸ���SZ���O�����k!_���-m�s�	Еⱒ�2��Z,F�l�@r��=!c� g"N�'YJ8����3�"e}�#(�hH��܄R9��}����l�g�5�8+����������#IS��#��^ ��]6Pmm7�")�c�+�+7CS�E�&���zJ�4Z���(�65�ǃ���_!��~�s/Z�䶃^9[SҐ�`�W"�(V̔�7�f8�U�
�ٗ%��X����m8���rr�9�w�v�TT|?u���\J�Dm3�e&�Q$=^ �/Qi�kJ�/z�.��(�n%�Z��3�I�\�/��9W����^��z��_�3��%ύ����.3��}T�,�F䠹u�S|,�\ÁRJ4���/8oogG��o�/qg ����	2�"��ɒ2���r�)0F{���gnV�Y���8��L��-:�����j;�
���UZ�He����7�/W-KI���iԬt=H$$&X��<��ߊup;K<P1���H�y0K���FH	A�([5M�F��6i�g�^w�Y�8 #0����_�BD����BL����)<���17��w+�Z����1����!��D�T�55�D�ri��³=��k�����A��$~0@9b��15�H	�T+�IoY����ՀپTO�48+f+[q �_��d�P���#1f���}���'�Ai�Ҵ�tS����PG�]ډ�9����[Ud-�E��s(��{�4x��@wovN��LE� jP*�i1���0���T4�C/�Q���D��_���aNiqH�� Y�[�\,��|�`3�l�Y��[�:]�/Ov�\0h����%b�v4\�%l�
C~~\����W�u�bQ�Q=˹D?�%�f5Qls�і|�����Ԙ������u�9%ҙB��qp�<g�1`1��~η�3������0:{�;�;����>j/, �*�:	�)HݼӅp�uC�D0�W��T���˪*�_���:E؎�Ev�Q�rd>��R�s��X�#�^�t+�Ϯ������~�M�'�
�Ʌ��C��$-�3�cƃ�|�h�*!��^]���.^{�;N�@�>�L�Aށ�MmHvQ�+���õK������͔��DmaO�n�nW3E�#C��
�0��9��h�8�մ�KR]�d�X�����2Cn�]��)����6�PТ�	���-B4Bʛ{�V�+9�9`bg=��Q�;J*���(Mw���ě5hV;��#����m�U��=;�4n�/r7�ю���Y�����O���DN����qZ�X�ˍ�H)�ߐ���a��Eu�G �v�W�;|@6�j���/�
��t�ka�����o���� ��t�4՘)_쑘�����t�
e������b�2��B$�X�<���<�~s#�7,xxҞU[�Ä��ozs�
�GM���9�V�l�kO�O�;���W'o�`*���.�����_a���С���Ulq�,1��6��s�҄��;$"���z�����{B��pȆ��Z���	��R �Zj��B�FM\��p�m���VnU�=��6���ڃ��޼�(a(�5��֪�d���XV�+<�ԃ�/�6�'x�p�E��`��y�	���/P�m�+�h@�?i���A��@x}YU��L�gV8!@K�`�|��:��yN�!NW�y�ɱ� ؋)�	�5w�&.�Ȋ�e��|gp�F��] K��Ɋ,�#l*��h����_���>�X~g�<Ѧ���Ak����k���6ň�xϵ��!|�f�x!��v��qk+^I�b@��������е���-��,�7lI�a�#��֭. N�{ex?�)B0������,��I�8E�C��D����9�����anA�}�R	��/��2z]����]-�~H����8�-ׇ�+���.�T��;n�jg����E��&�N�0�_���6��������r��.��͍���(~� ��N_��݈!��n�=`j
X��������[�GO]Y��#'O;$y�N(�q�I׵��s3c��o���6�j0Q�e_z%}��(qѰ�U�p8
�c�1R���N�c��?e�m��	�H�2�]�\2ht�{=BN�0Eޣ�����gh��i?���>�J�'�y�1��r�_�E>��1u��2�;2k",�	���p.NDNl�T8�_�9>j9�h�����K����E�+_�� �ey����O��]�i�htDJ?Π��J�r=ד�
 w'*��%�	I�g�	��BX�2>܂0�Pfl�'�8R1��%&���H8�� .G�Q�J��jp�x�'f��|�:�G�^�6�c<�1[�B:�I�;�(Ja�W����Hܩ\Bb��[M�d6�s�6��G2S�,Fw�sO[�:��5h��k^O/?m�b*"iK*�gڧ��t���ax�pr���$��]�6��i�։�Y0�ī$jسZ���R@�]�LO����L�!'B�f 1�'�iz�j�}�Nϡ%f��m}N�F�.�>$F*�0�M�'��}l����*Y�*AЙ	�^�̷�M����9��x�'Fu�>R6��~	��͡̈́Vݧ�\�/o�!�Aj4[v�fpH].��	8ׯ+��+���3Ϭ��ہ���W��8��)���D=�=�=pÆ� ��bGzZL���H\3US(�}D'Wx����6�����&����^�����.����y�]�3dMAF�ۀ�L�(_@Yx��5�8?�`�e��A��k���0JG��v�^���%�*�c��2C_�UN֭KI��_��Ge�BU/9ȅ����� �@J}�l�Ns��}�BtZ{�\~,D#!�`�ɑ��o��5J�pi}��x���Џ�yc�>&��2.�q�m��5����Q����S9ۖo�dٴa����|a;1�W��I0(��wo8�HV^����9ۡy�������}�����#(��/Œp+?[�(IBL�-%V�b�9n��#��Y�/8E{aV�;�0����ϱ(84q)l���BO.��B&�֩G �gĄ�����E�Bꃁg֌�*�?��
X�YN~O������t^��&��+ˍ�!�$��[`�ۈf��N��SI�9�n	����KB��hmg�B���Z��T�Ζ��g)�"[�FD���q����um���Z��BVE��NaF����<Z�6�أ��y_�#�P��h.5��I�v�V��0�gjp5H���7�S�y�4�DQ�PP?�S�R�3	(Q<7��,��r���
ss�t�����m��^���xGw�V��K�WïNi�i�x Iߚ�&��4&�V[KU%��e�!����v�IFJ�!��'�CSԊ��5a�ʸ۰_���
�+|j����n�FT% �͔�Vԏ��yee����k!�qG�~Ʋ�y��i���j�m՚nC��<	v�R�w:�l��a���M��{�Tf���嵬�܏سՍR0���7[���%uEX�8���j'P��c��G�*i�/2�EX��w.m�t.�T���6p)��Vb��&۰%��xyl�%tP:b̈́��Ĳ�	����ȹ.�4ސ��Op��[uɆ�������Z'���u�8ח���_�cM~a���Y/xq7�����u�'��w�_��Y+��hu�_'+I��e�trM F���̅�D��to>dUõ��R)=cG�2�6w��!#��cU�����p�_��О_U�B�E'�s�dUi���d0��7���ʮ��N��,Vo�GԙG9WaN�-rs��_��K�8 �Iv�/���g\Ġ�Jv�^���5N��Vp);`�=���W�ɿ����kO՘�[��0���T��m�m*�T���f��FӀi�����>� !���^̝R��A�rF���^_	2r�V� p��q-WxbGoC��Hg�SЦ+N��^���#��d&�lO�+������SC]!�*�~���M�y9S�LU]�5�����R��+��F���c��������J���/�~=�FR���h��c���f.K?4�<�qf H��UQ�ݾ��mWy�8�kÆ� djm��#���|NJ�,��G�\N��G��C�3�'�[9��r���`�]��[ڔ�}�g��]����>:q{Y�;�J