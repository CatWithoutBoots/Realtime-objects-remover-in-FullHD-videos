��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&r�F���oh���t����v���@�i]wpPA�Sf��dG�G�����$f�?�yi����lmU<�9c	N��O��\VJ�!��Xzа"��Pƫ-�ۇ)_1�w���E�$����4�]�8B�j��(Ɖ�V��iK���y�'��B���r��W�,A�Ιs'��$���p�^S:��%pS��A[c=�=�\8�&��R�<�h�p��u��C�����aq������JɼP�tE���Y��)0&�"�F�,�ȃ�t-{��Q	�����p)V���oJ��}N}�c���pQ�}7b5�E)���H��W����P#>�|f=#��k�7�!]��x�kRL�7Aý7v)0y�K:��[�j5���S_��Q#V;;^Gm�CbO��ߧ����E)o �]�z���K k��~�h_��n|�E�"��k;�O C��ݮ]���og� �j��*���p����w���e2F�d�&�,� JEނ|��
#���y���J��������kщ�^�J@�2N��S3�~��Z��9�y��MC���-Y[G"����H����Fiƅ[;QWj�2:O��N�&�qF)?�G��S����x4+i�D�*��f�$rmG�\�[�V9	d
}A�G�S�9�Q��b�J��s��2�2�u�O]�O^� �f�xs�+)<wd����Ƹ� n�j`!��a+��������!��Ӳ�Sk�7�4\�P$��(�E�3wv�;�W�a/Z5�^��b{@��<�d�4+-���;3�@��i�Xn� V��ʜҰ�	��7N���1���(�}y�ӫ�L�"�e��K�6؆*Ur�� �w��$Be5Q�9�f#~������u	�J�%�+��?�Uo�|��b䙙��ͅ��c��'�e.�kU��iX��,)nɗ;F����%�E�s�f�ĩh�F9���sףIs6���7E��(Q_��K�jT��˼�n-]�3V*�BX�c6��7�A_/��7�����4N|��w\��ĳ�".[>�U,3W�s�k���AτT�z:#qC"%���l�/�4���������8/���\��	bm��xW���X�T�߭u��bt�nN��26A��?q�J���2|k�ֳ���1ć/P��'�!e�]TޝP�NdtQ��+��y�w�������/��l�5����tд���ۘ�X��^'���:��w8���T�U�DH�!,� �������*��6�R�a-���]�z]4�s����n�����M�OZğ��*��� �p��Τ=�n��f0�r�2��EY�oG�,mGM$v=���%��c��Ѯd�o�&��!Y�8�[І�<�a�?������'��eN�s�T���ę�3�n�Ki;�*��K+��Y�e���l��I*7$a.�U�������y�dq�a<�EЋ���(�����Ї�i5I�^�Xu�f5=dF�%D��6"Z~�dx�:TA$q@%X]�~p�fz��E��F+l���ED���G7JU�7���o�M������3	��=;���0�_�t���,7��G��ɭ������C��hDwL�
cY����Z�C�s��j+���ض������n�AHˠ�l�S���7pN��γ��.��Op�8h-#�h�����#��%�~�c'��A�q�Q2d[�?5���M��ji���On�Pq�(�(]_R��kQۺpX)̴���%aQ��s�=M�@(���q+R��'DH3��rw�W폞�ƫ��`�������^������ֵ���'�tQt���8 =���{Zķli��vA$��$����r��m����M�E�M|jڲ�=��	�c� ����)��VB�o�b^)�z�ΤұC��+m��: ^��O!!>���c��A�wJ��&*#�C`϶uVY<4/?rIQYm�.��k}����:�������5a`6!�]����RFŇ��SK������C��g5�$0XUb��� >A)L:o����f�Fy�Ȣ�E�x�k�f��U��+�ca�L��m �[T���z��Ɓ���6Q$-{�9<A��G��AM�jG*����D �{������kϑm���0�ˇ��2���8��dC9�`����`��&��,@�MO���}���W6��-�/��{�QH�,虅gas��Oe4���K#9�]w�*=��6�|��@e�N���W��fY���[B��<+Y�1�������aK�K�R@č�Q7�Ѩ�f�_y;tm@,P�����@Y�-�ǷhH+ ����성^��=�;��sV;=v��j��)Е����N��S���H?���L��v/*�hμ�\r�x��N�<��Տ� 1G�E=+Yuʸ5��G=$?���,!����M}��ې4�\S��;�`�5jY^��};���(p�;}��?rĐ���˳>
铉��A+!٣�k��ω�x�*.�vNm��� �l�(?����\�{�ڽ�1��m{u� �ZS���+e��n�w�\8�M��r�*{/���Z MJH	y�0AR���0�>hsWH�� IF�I������s��0|m(�q$<���+�W������T!�~�c��wv3l��Ԭ�>��ˢ�����������S��J���ױ�n�������-;v}�Bg�kLyeE�'��H�,R�?���y�Y�&"�ش�aW�Guʨ�=��j*�	dXӉ:�n�D�p����Q��ϕʣ��U�q�z�3M.&b������:\�@Ǵ�\�䆞�7+�$���Q\�4�� �G�S7r�k�^��r�:~ ��Wz�:h(��!񅆊�[�>=}Θ���Rk����g#W�s�l&��.����)Ii:�GI&�M\ʸ��ܼ9UP���jB�� ��##�[�A1�֊����I�kcZ��!w�r4
+]�����0����	6%�Ffߏ�M_����<t�<2��z>�w��zW�e�¯n�; ͩȒ��\m�&םv��~?nV��'��T��M��Mv��~��b94���]���F�;�c�J����<#Ŋ"=y�:��9;No/`��	��x���;�*��!,����b�N�mK�K���:>n��ՁV���ܞ�@�����A����1F�?w:u�8F�Z���p����D&�&�Vt���^y�|�"���}����n�C*k��}7�A>f���Vٓ�H�T���+�۫:��oRQT�Io�^��K8$:���(0�h����s��0B��wm����BRP���}����f��.�aZ���M��$��5��nU���v4rq,��ۢ$H&|'�󶦮�!E�X��ȴ���� #gl8HL{�~t��ѕ`lY^r~֨[�����NC�<Z٢]�d�rM'j�.|��Tp��M�N��h�l� Z� ��� ���? (��R����y�O8��n������OK�������2z{�l-�y�?��~��ȅ��<�	������e�@����뽆�}��Q���*T/r{b�_'h,!/_���c���ɕmY��+��h���#�O���o�9#�^�=/?�,O�h1��`]�p�3�c�*�ۏtjy�-��xx��4���0DW&�p
"YlBpv��¦K����jK�-�y�0������^v/TMV����V��vd�f�3�)�(lj!�Q����0.ɓ�.4�API��2�@�&�sT����\��sb�}�l��Ur[��ŷ�������[���q#���3v�7�.`���+���d�]g8Gz�.��%r��nӋ���iA�4��c~7�uᩨ�=�M��KDDv��<V�!:J���4�5S[G:pbڇپ���%�kA�'5�쀠ɰ�FȒl:+�阣Z3��<����50 |t:��M����"/�-܄��|=��Ǆx|�R����ZCQ�C�l������.y'Y���:��
;�}�j�����̈��+������"��8��J�%-�A�K'Q�h�@�xU� ^	�d��wȮ�R3;��Y��4���f��r�W3�����|#x�����L!�Ȋ�>P� �z��'���g�jW�'�!����e#Q����I�KX2nj�U�L��V<�ؾV<�v`�k�_^�"\+�`LH���,o�I����`�?�=9�".��?�K����C��l���y���i�� �T�VBZ��~A�S_Xh���ׄ�����B~��z�`�eI��L >ں|hc�cS0���/�tR�+Έ���`�p�fչ�p��Z@�����!�~{�O�b9P.�Rg(l��Q0�Z��j�GxΆex$����4���E��-��ہ���!˲xJW�r�Ya�/�6�TB�}ꖵ�*�9f�f�o��bZ���/ϛ������E�������������B�.Bvƍ;�r�Ͱ�Ab0�kuz-�ҏ�E{?y�%>u)���� �T�RJ��^����/)�L�A��l�X��sE/E.;�M-Ny����,<{B���@��+,"R� )aɆc�i(:)F�##d�R��OV��l�|�׫�!�TV��f5|˟T�<;�JD̄��I�z�A>j����!����4W���U"��(%�}.`���}�*s����m�/�]��D�G�/�Ii�SНv���`��p�6	l������gOnl(��-,�֏����-2Y��`�_�=��?��]PY�,<�4�,�x?A�f����GL�(��5�5*{'|`����!S��f�/���J����瀜����L"����;�S���5�"�pO���c̩���pP���3A��u�cM����.�8s�='��h�o*>�`���o&#h�hejvj3tL`2�+Laa�e��3��#�F.���$9(H78z�U`]�$���ǁ����Ah?V���m��q��ӗ����L�ãJ�c)C)F=W�� ��Uɪ�bz����(I{�6�q�'�D�"��g���j���I��w�ݬ����l��1&��	}���9�.bx�>�L��<�!%[�F��9�{6�\�P� ���X�d�����^�^��M(�_�W$�6+a�Ι1Bkf-^I_~,�7���Ȗn{2�5�������0�Z_�#Cr���I6<Ѷ�_K����,�"�#N�=����YO�K%������:�!�i�Վ�9i�ç���e�XSBy*�J��c��9��J��&�BJ��	k���z�|ZiL�K����Ɍ���D�2���^��`β��	�
�%]GNI��(Ǜ��}G��{���s]5!��&��q�y{9n��ϫ1FG:��4���{�2V/-�4�
�6��v�f�z-�v�Ș�H���2ڀ�"��]���rܠ����P�A|�5�r�Gx7 <�q��N��������"���r��'V7�}�eФ�؈?H���,X݄�l6�ȩ6�q7�'�G�z+t��*>�sy&D��ږe�*�Б�y�:�iI���4=���Q�O�N���rI��G���P�Y��є�=1�,�&�9��o�u���+�tz���a���Z�k�"LLk��x�l����$��|�T�<i4���B-0��+M���F�bcg~�>��H��_m?�r�	N�u4�<�-D����9{=���u��M��6� �e@;���ԙ�����wo�$G���"��&է+q�4��#a�	TSy�3�FBY�Y%�Ӈ��8pӐ���\����-����}ިH��C��mB
�1
_=M"�#�pD�-�_Q�6'��E�_u��돇���B����0���P.�,&��X~��T�����8 "*p ���G����'�O���UQK��2�?Fz�����~e$��I%�+չ�nY���/�{#�Xi�&Qb�,R	�S2��3B��zx�6j�{F꒴ӵ/E�@�t�p�/�+YZ�ˇ��g��z�+�T�l�mk�S!�4�P3��wx���q(k�
���p��iB9iΌ��+	HZ��3�eQO�Wm���w
=���Ktfx��[X��M��K�!n���%7�r�Û����.��l��i�v\�I0�;8�A<���"�����Y ��A�^�Gs�◔�k�V�%`H:ME]���/�k��C�2Ϻ�ж2[��$�:-�(��~~N�U�!����%)���p��Fb \Y�'��b��(��V���Ǎm�Q�bZٟ��y3f&f��B��!�����Bm��f�����5�+��3���������Y2S�
�n�4Պû���⺹��o��uo�����@�o�1����'G���}vGq�<0����dt��o�*�H�H���`3H	�'/q�FW�-�@u/�c��s`��O:�S�2RlV���"89j)��?���&Ǚ]s֒���Tl����y1Xt[�������8
�_�VM���gt����.(������0��iF�� �uf=��USǬt���7�&�I�h�h��I
CKm�3Xz�Ҟ�g>k�	I���Xc&�NՒJdU�b�ƈ�rV�4�����-Fv�R�@8��,���˲����*��H������"�0�Yx!�"�O�ePo�*;��6�j�>@u�'(�2�t��9�nÌ�G�0�|k�k������� f��vJ�.�k���ŏ�n��r�'�nN������X�ք�^�ހ���ϝ�{%�8(�+�K;����+�r�[p�lv���_-	�΅�P3/�=��s;��d��<���!=5��%�s=��>+mƃ����aE�7I��9�mp!�?Q��B�g�OX����n~���U�i�_�%��b�cbR(�q�#-��[q�o���Q��e;���8[��+)�
�*~A���������6h�]ٙ}��]�AfMZ��5���y��vHIt���+[G�NV���җ[ߣo7����^�~�p[���>�0i�G~p`���B��o�;z�Q$�+f���+�0�@e�J��
qVf�xވ�T���>F��6|�8A��فT���2��7%���Xa�x�Kj�������U΂�->
�ډ�Ԡ�KȺc��TP ���i}Ļ
�2 kd�㪸���j���!tN;���%Q@�y'��z�gOE3�`�R���"9;�ޝT1�6��,2��n��HAt��o[d`1�s1�4�7�p�:a��ƺ�B���)f�i?O���.*��yx��#�`�Pw�V��	�w����y�Ǧ��vJ'��<�v��d�i��X��Ў(UH����4��sn�J���q�/.
������G�!ݑ,y�7����ex�8A�� n�D��٫
>n<?J:��%� �b�� �ՆB�3j���lĭ2j�ni�.� J%�}�i;A�<�(�����Ӥ7ܴ�:��;i�|t� "b�A5�<�P6*��6ea䛄/��}Q�Ɲm�2UАXKt�J�	q·���W���[�e�v��nY�(Р3f�7�=*K�����4��4�E���
�����=�j��;�t�:w#���,Λ�2"�OS�[����[{�Դ$1�3"g�wE%����,x1���X j�H�y�:\�bR�����S<43?����فt ƵM��ñQ�t�l�v�or�P����UGv>1z��ʽޫ"/��r�-M�z~���Kx<����n�������I�bX�&Ʌ�j�W2<h�;��Px;�v{+��X)���0*��h�\B��!w��H���b�%���-�C�[��W��锊��w�I���������u����x�)V�]E2$�؅�!'�K�)���u3E
W�؞~?`7�MX3�V�F�m ���u5������y=ܰx�z�C��77r̤���ࠡ�S�ޯ��`�����Q���>�o
+71����Mz:ʶ��c]��4���zL��2�������0?t��4�d���44f���\��
����V~0���Q:΀��Y��,���c:%%��i���D�9�f�^�T�E�T
yf6�M&�b�܅G ��v'�3'n�r�&�+'�l=L]<�&�%��ot]<&Ka��L�wf��C�5�� '{��yTn����`�\��5�2����k�GP�J��zg��U�0F7UUf΋�}��@i;��+�j���[��D�-.9+�v��'��[���Z�,�X��*�A8E��\��SD�'�� �6�X�j�"mn����R�n撀\�No�
"�b ��l�M�)Ƶ�~��&�G*>��ܳG����E��n1���n���e��������w�ɍ��!q�Ϥ�{�����*D�9ad��企�Ǻ�U-S��Gκ��+��t|Qu�U��)���N5*�b�d���B}xm��ζoe��崀E��2V`i��xT�1f�H����l@R�~�����!e���8��w�^A�9�(#�G��n��n	�D�K�aW�(�^��'=�G�ʡR���