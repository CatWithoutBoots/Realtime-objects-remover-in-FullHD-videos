��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&r�F���oh��7�K=U�u�X���eת����N��/��Wc�4��@Ĕ����,||<c¤p'k��ė�{�%1�-�-_��J6�-�#dV>������������r�
O#ENM�	.Na_��	��x�r�N"Ȩ-ëVj�#9c��l[�����l�i��g�C��K6�9:�Uu{���A��
�(nBU�����z��h��f�P�P_�;��#�S�P�i��A��5sx�!��ĜX����+ʂ��g�?J�4]�kY������?B9�T(��oo���;L�Ļ�B<!%UAB��PW1|E�N�m+��l�* *J����5V�Nkdx�	𫷰%I��X\H�o- �h�yi<6�["t!�#�wLK���G�zc��{�^ҽ&�bOU\����J�I��^t� �X��
���Ӕ�['�/\L ���$��ۣ#ZK&2M��
~�u��^o� �af�u���(�O�� �P�n������缿=��ɉθ̓��ʭ(�A�,{��;�(е�t2�,����"ۼ�����l�L1bи(̡"^ ���� Y�ǌ�q�����<_�'������'�{��7�z�OU(���G �洼eaa�2b���ܲ�z�y����}�V���V@�fG�ע��K	0r�n�v�#|W�K���?�7{NS6�_�v�mӛ�]I�»��I��[,��:Eăs�yܴ�aqG5���������惽>'!y�Aģ��T�仢��A�98e�e~�pdY\�� ��Unп�=�m���]0ĝ53�1p�ODJ���
� s0�eZ�%����ke��7�#P"��ܖJJiY�<�h��شMb�+�4|n*?c�B�u�%��s�n����Z��
H��hx٘+���$/�#�D>�����U̹z����gV,�T!�N�U��������a�"V�\�ź�b�-J�y������D��ᩖL���&�rG�S�W�x�Z&,gSU��N���	v=���c�T�F�)J��6����k��R��p�$��=A���o�c�xMrId�Kg�b�e���r�[���䫈H�?k�)����,��=03�R&�oP�D��"�i��^:@p��yD��95�i�#0mK]&R�v�i>XW�;`�.>G�;�ʟ���2�d���B�`6=�S٩Іq�ܖJ�Jߺ0�M��c�яFYӣ�v�3�c��}����v��D�%�w��,���Fu�H{�����f2_���>(�V���8�.�&+��e�z�M��.��g�Urf+@��ۄvV�BG QZ���6����W6#�_,v����Ѻ�x�m�}օ_�> 	����a�gWE��"n�����LL�V-��«�IN��m��r�4���|��]C-�Z��d7������ҡV�Cr ַ8-1�ɥ0E��)�Ƕ_p$��;�HG�
��E�3vB��w5F
k���뾚I-�0�vWl�?XE�A�.���1���1��x�:"���X��� �%m�&2=��P����m�^i���-��>�];��p\騽�{�7��@��C~$ή<UY<�:e]�ݲ#R��Չ�\e���}��xO�"��/!�N���gN�+J��dN���fN�QT�w���I�v]D�»9.y�z����I*:B&�O��JG-��y�!�!�������/��-w!��|��u�W���FZ�D-�_�f�r%��G��<��`nm��a�� �	:?��<���rxѼ�>:�vH�Lo�΀q����*"%9�@yZ`�u�a'o�,�Ǐ�5�e�>����&�M��길=	��:�5IL�J������E�� �_�tK����I1���$e�wg�#4�GagB�n�8�M'�+&R��>�pwzN�,�\P�Tg�7�~^�z�&)�
�m{ST��w�q��4�X���CU�*\}�g$�M*��35��B;^X])H�h��?��|��w�$Osy�𾚾F+�8�ױ���{��X��Y��c�$|(�?~�`w�͸ȥ���7��9�P�>�Ȩ� -�`�ig� F؉���Ց�g�%ru������<_��Ot^L-���J��R��~�@Q�%ّ/J�