��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&��^L�h�m��uXҰW�J�G��!���9ǹ�U3}���|	V��r>a��pZ"M����SK�����Ł�G�8�Ek��;v�F7-�̏뽅/��C<V�Ar� ��FE��u��k?����u��S�/��|7|�P>� /d�����#�H�,�?�V���*̟ő����t�ҫ���O��0��(T���,jAE :���J��Җ�������j���զ	��<"�ф�x�^ll}DB�+d�0�$m� �O�Jkz�Fy7 u���+����|Tg�Q:N$[������l/��R�������'�|�ٳ'��RW��vƙjgl����������j��l�^�1�^��q��o�����ut��)����ì�˝�����L	v��;֜��)�ٸ��n��5��'&�Ƌ���2y5��O�����V���k:+��#��V�&���e�څ�]��4�������A{Q�&X��G�ovq�p��/�F�� Bլü��{?�wF�U�$j��~����K�P%�M:�?~7�fvс��&������t�0H���S_Wj��Ln^���룧_��)�@�trR_n.��=8��Q-X�`�w� h���0~N���F|;���>ۍO� �0�k�8���߮ɒG�s�\
<M�����캬R���B�T�-X(c�)#-��Y����=E$67��u"�R��ɍE�+g̊�t�o�eݴ���hzO����b��8�e��"Quz�Rw���?p)P�a~�����"��T#^h/��٪�|ӄ��䔁\�g��IiYG�v^�U�%��V�*!���t��f���tgݿ㮭���hww/92Z�pcSN�>�E0�������$�ә;H%T��A��U��v*}"�O�DS��o7^Z?�61�{Q�� ���(�Ix�wH���\�0���k��D����ѯNH.y�T�m��"$�x�\ �"�M�Փe^�C�E4�E�MW��[�h�Ox��z ���Z�ΰ`��%��s�98E�6���P��v�N���R��G<^>��g^1�;���Z��,&���"���i5�G��3@am�ߪ����\+�@_6XZA,�GP񐦜Ⱦs)��I�1Z��'3	�P���)��(�
��r��	p�2o#�ST�9A�������/�zn~�$���Qf���T�IL�Fh��O��[�ƙ����$C�w�d,�12�ΐ0��W�7#��)��F�����o����R�s�7��
TumW>���M� ����:Ṓb�o6��FL����NC���J�U9N��9 %4���]p�1 �L�!�ڝ��(r=ŋ(��tu�V=�̓���o�y�'"qV�C���ܥ�%���`I��X���н*����b�~�J���C&?80eF6�.�H���h+�������0;�о4S��/F���0BcY�(.�X<��JP4D4�uR�S	�Q�k=sj
�����nP���j݈/�X��&�|��ɚ9Z��C��@��}�N�͇�$���d�>e��O����U���{�x��zV�
6b6p��f�|��k����
x�dT��F�9QJ�zINZ.y/'����abQY�j:�LOzt\P������(Y��i�p��A�X;�`�P���m��Ǣ�l�}�d��U	~�y��h��xt��5g��j��L0��Е=z\5��V�t�_�m�.��{�/�U��$��fؤ�1Btsd�>�6:q�*��0�Ϙ��=�| }h�G /�c�&<;�'a#����s� q�`�[\�,�y�h���e�ϣ��Q~�ԖFϣ�d@�+�$_=�,��莙۰������/��.�{�����ۡ���}hDF�bG�պ�4+���ڪ�p�(V��`�UE�����d{�f�wI�@�[>G�O	�'H�	�`���Sւ��40j�Ѧ� I�z�@Ϩ�Oh�G!t��[���q��%z�������s��8 U�U�D����wO��6��$�g��"�d�>X����`��bzYmR�o=!�N�Z��I��\>�ft�l�޷��r�'���9cr8����-r��ڢ/���`WiI��=�r����V�(�� '�����o����ӅEK{� -���O��7}o�,��Õ?��%��Ʌ� Uы9��*����!�7�N���\�R�I2�;Wl7����a�{�B����7�߼�W�]~��!����@Gн�(E	꾞����n��L͝�/�?���d#x�� rH8����*���%�Zh�`�8�4���I����`B Fs�=���yC��0CCع]�/��(�߲�]�h���)�]�A����C��V�(>�|(8�/Ñ�
��槟Da�|��Yq�[�X�@����fQ�)����=9X�_�y=I��߾h�vs���R�����B�ɟ�d����-�tY� ��q��W{#.�صrU�`���~0�e`�vT4��
�N���A�L�o��}n����tp��td:t� ���}�6p��'�j��ALي�D1���(�l�L�.&S92�ߣ�G	��co��O��r�&��Bc^��|^�p��]�qX�T��� �Ky/\h����@��vC�.����3m�;��G�O�f��+2@G#����&Z{cF����5(Ջ�M�����˲F"g���IT�Q!\�-�c-�77�7��ەР�Đ��U���2��5��-3�I�-���<��W#��"}�=SR�,V��t9�vDZX���	�G{��Κ��r;k*���J��v5|�NY�|���>�ڔ1_�ۅ%;����E/�����D�_�Nv�E��.G/�*�Nt(��	t-�<�o��>�� }��	����PK���D4E���+�xi�9�1�Ok��������O#�� �aI�Z����x�Oo�f=Kް5���R/k�W�$�5x9���o1���^;� ������)�UӅ�T��f,<��Ͳ�P;�;J�BÌ�uoYi$��sWd�LC�9�sH�	��7�Ao V1o�2���t���^����?X���������L���q�t��[�˺�j�Ίz�,��Q	����cY��i#��#�*�G6b�֕�lE�PP|vQ��Uӗ�T�9rŗS�B��=(H�+�|�/�9��RRa��k���rh���		��x�%��PPk������6�_&0"z^O
ܗ FA�*ͅ��릸S�_�ȾW���U�s7�gO|���cl|/C��O��],}�����M>D��"��#�lי�
&�y�BZ�f�/�6&yN�����G� ���X&���P���j�3��n�P؁�Y�k�e�UN�sm�%�� ����fd[�,0p��侲�jM[D<{�&�4��c���F�Q�We�Ά{G�
o��F���f��D�{���%o�2D�QKd���@� �]�Y5Z.�� ���R)m�l5��-���&����h8f!�Գ8X �?���fy#��L��ױv��Ӓ	$�a.�>Z�|�?��`��/F3b��lO�
rI� ��L
Bp���h}���X��u�+]�eg�υ���U��X��OAN<E���-	��z/���n>��=�������� C�����U�����D����r��r���֑��ݷ��
E��Gsm ��~��Z��O�%�wp_[J�g���K�ðS�?4G���ѮϘ8�u�=9͐lY��+��|f!֩X�c�M�O& `�__>��k8�%fK����
,��%j9ߗj��bX�\����г���n]��3�^~yĲ�O��S��W�l��6�8�0�e�>�R ��Q��<��BJO^]-��@g�W��C���|���z��I ���?qq�"��?&���ۮH�����0b���D�K��T$8}�=��:�3�.����{dI�ˑ����\����_�| l�ijB���.W,�!y�K4FS�	i��D���-�������ՊC9��m����=�_�IS w����j�ɔZ#l�.:�FA�ue<���ɿ�|yj��&�[��\t�qu+|P�廲����Ys�NZTp'��)Z�S��>n�k�ysdy�n�.��/"��7�AF���J}�v\�vbO����(l�c���z��N���_�W'�,	�L$���K������ʋ��@Q�-n�����U,��f��o5}RS���4���3�������1������z���i��wbm%������`����D
�,��;4~��3<]�q���[�踱�C�����I�/C^ıa���	%R�.lˢ�A�qDfF�9�e�"2�If޾xȶ�jS/}a�G���ި�T�S'�����:%���0�&ϔ�dյ+Y��wk�y�|�֭(���^��4Gn,�>�Є,�D�!�'�n4�`�/����Ć��َ=�� ������d��u}�(���J�"���K��O�Ea��]��Ѓ]Z����U<�Q��H��@�>h%�g���B~�D��(�JY$���2;
NQ��/fs���l��~+U���S����UO��0��n|�YT����Ѷ-��Y�-�H���e��Pۯ���v�b����SK �@ ��b4M/a���4>N|�Wa#��%��ƿ@��|e���&w[bGc��8(B��6�曂�\�x�
�e�$��;�ϔ�,��Q�U��dTe`ȉK�A|�0�M �xL0<3@�d�N��ki�b�	*�����S�R"���a���W�6M0'ڇ����-�� _Z�[GDM!�gEC���IFH���\�Vð�[�x�ĭ���c�c�u�?�噺���%QL��D҂`�.��:ʯ�1\�eI ��a���^�0��͛h��s�օ�榪��H�F$�	6K��0�n"�M��K�W����y�Om)��r�9p�B�����?�ca�u��<ڋ��V�V'��G�?�Y&�K����;����8e�z	�:�\ 5��lߢs����Qƥ?��i��3H�
��F�Gn�B�Ś+��Ԧ^���RR�ׯ{�:���n�����)�'/�"�b���em� KY�*EM<\|�/�ӀI��x�9h��[u,J�V�,�Mm̡�(=�M�p%Y��L�wJN$��q��kk8�F��n}�R�����tW` "lN����=��~��I ��09�y&$�Z�M�8����l}��k<�d���?/p� G�2�V��kԺ�w�X�y]X��.��	m//�uQhC��7T_�����9�������D�-�	��%�~��>�D��ż�=���N��%^�����uق4.�l�'ש֣G%-�a-��b o�?�m���E�A/��`��5�Lo�;+��,Gn&��6�'����׻6�E����
|����ً]�Y�O�}#�m�YF���uL�}7�T�],$ѧꅡ�Ҍ[�����Դ��{�a�c��c�ٟ��<؂߇_ �S6���a�l�Uh��ת%!�#��Cʏ�&�.��