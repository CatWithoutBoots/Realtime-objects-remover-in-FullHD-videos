��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&��^L�h�m��uXҰ<.`D�iL[u%y��2�T��ͪt��R7��b:t������g(p4�b�U$! C��bas����>D�����`�ڌ�ܴ�kt���o�A��Wް�CY��?�h���m�j�C��6�:�s�ghz����rgVL����G��N�=���FP��Ӷ:�s>���J�Zʅ�ۇvaA�}o�;�*@h�M���_�~*tf����J��U+_
w2��4����J>��1ɇg�@+si�VlX�&Sg��;�͂�.�6�nh���N�>�S��0���N��kDWCR��Q@3�EXR�QRтx0Լپ��%OdKc�DP��p��Y���0U�+�*��oJr/#{�~�^����NPB�⋇�,Kl+7�X�ۼ�z��K�7��bXh�SFeJ��$����UT�r=���.x\n�Y�t��E���o$x\�{n�9�VH/���k,VjR��fM�-o�G/�[b���Xh�I ��\o��=�+�k�˒˽�ݨ�TE��:w�������	X\���z�F=�i��>���D��C��F?�sſj��	=��]N���Ol��5{�.���U�p��(��KA�O+�t(��Ƒz��DFi9�i��S j��]�T���@��a@��&�Zq[�ӣ�^x��f7ò)wr���\К��ļ����&�+�Y�*�8���y��DH�Y,۪��Ә�+��*m
�J�ڽ�Z�L��o�{M�Q�# ]�W,���Z<�_)N�]0�J�H*x�-t��Ph@� "Jd:���+qT�}�������'O����}u+���`��z�Xs�=��
��h�C���>��]P�~��n�Z8y 6��N	���=/�KU�A2��,\ �ʰ�yȣ
�c�nhW{]%#���k��P��֐�r�.�l�d� m[��S���z��I�����{�zk�r�׌$���s�4�P���6`�s��7�|/j|��}}&�� �̻�Q+z�j.��lI_�8
l�<A��4Ӕ77a
2��닮�h{���r��7�AM��o'\��|"I3�����>�_ ӷ��e��D���O����ǹ�~P��E�݋�d8��eɼɠF����F��H@������
��5������Xeb�c��a�u5�7o��H:��J�:��D��r��u�َ�n���#�[�$I�(F��nB���N������/O�v�@߁Ϝ�~+͹U�s�0�ϱ i*Ͳ�D����/�K����y߱)�)���-�8`՞e�ȋ�
�7��7%�ͧM$�%�����4`��7U(! �&u��{�ׄ!ZeH5:�u��:��&�b2t�Q	ݒ��$��ۂ�t� �N��<5#�^
�5—!NZ�A�r���47�Ah�Rr�����{|J?��b���� �����D�$�LT7�����<j_��v���.�FO敌�"����r���&���l��RY�<ă>Y�l�o0KAta��//og�}:;����͌v�
����ผ��ȗ��d�IhbrgWg{�a�듣/��b�̕�{ْh��F�v� 1��yЖG�JK[@$|�ǢU����pRp��*Ы��B�O"��5�S���L��K\��Rv৯��zKնb��m�a���_]!�ߌ�V�f}�P�)��aBI5Q�"�?=�y��;�Lt�vvB@o�U�7|ƙ�R��M��Q\�|�B7Y"�(��6ac���S�_U�^I1�g����ȶh�d,�'♈�*\@9B�l5�)4�����S(�թ��~����x��a����5��s�GCrC_�S�R�i+��˖)_x��%�6rL�J��������yX�v���p������#�2#.o�����m;FbG�x@D�lyh��U��/D�2GB͇��̌zx%�����[S,fk�fN�-6��.�@��۪�)}y��~<��N��H��"���/(wRb&�?�!�pʪ#;V_|�2m�ihקO1��]sEˈ�huƾ0���0~��E�g2��.c�f��y��&��&X����}u�	�x�c���ib�<{�Ø��9��B��@�B�[@I	_*����	ըk�)!Q|�p ���ƃ���j>& �_;�>x��P�O���t�(H�Bv�ڞgT��v�0���{fFѪ�6�̝\�,G��Tp$r�}�~q�Xk����Ӫ�x�j�i��-b������mP�'bF�����Z��>�[D�I (��"���O�y[�_4�r�*"ͭ���0����~{��\N*�5޽?N��b)�����\�C6r��ޛE�����\�!�	z�T z4�ܤ��`�4�֢r�j@O�� �g�����/�>w��d,���yė%֯��V�X��"٪?�ۓτ���� �b�G�R%�Q0���Q-����2$?�K.Dhq�G�У�{5�?�1�8Dy>�"r����?�E�I���3�C@܍�`G {1�J>;U.�8N��3�-��.`ӯ��8U��*�FA`�+�������q T�q���7S{
���1C�^���G��r�s^�-�b�r��8M��;��~c�q��I!� �] ]�2.��^i�q^ۻ��S��j������s�����x�F�CZ� ���k�	o� ��6��`=#��d&j2ϑ���Ͼ�򇩟��ZY?`ե��ٞ"t��Dq�k56  H�s�_�r�Ę=�̻I  �g��9���㘗��	uHWEԩѡgu�4�U/V���Yy
y���u�ln&]5�E}h}+|�x/�E��b�!MV݊M���^ڝ�<���v#��#@BgO��OW��'�,��4w�HKNi��g�4�Np�&b��  ��j�\�85�%�bt��F��aM��[l�RF��'�_߫'H�x5!���
�7�r3�"��ˊ��Y��WLH��&.��hksǚN���闾��� �������_6�ж�:U���Y�7���sR��M�'P�ɬ���U>�8+J��o�N�H��@��
���.@�k g�aa����)��1]@OQ
���]_W��[�6{m���C�ZE�o��m3\su��"}�G��V/]�Y�������~D��&q#�D7���>%��!0ﰼU����]Õ"0�e$,>Ԏg��Ǥ�C�	���?�`��ル�M�]�Ο߯a��W*�mH�t���1�p�ǰ�-�g<{�P4�Y6�f-.5J��
��Xd~�TNk̉�
��EqY[�A;�l�v�P��c�f�P�>��`ګ���W��M>��а� ��Y<�B��E���#��Q�h�k:�qf�Ka�m:�ob&H�pio�[����+d������A������V�����M��]�������3�Tj�7����5_ҭy��r�mX��n�+7�8�d��k�țX���;�����HG<^�Fo�9v�eU���a�!W\UOH�����	������� �.%�����fLUh���;Vu>�� �7G);u���q0Hh��*�
�F���0
�f[�_k�P�1��8c�L�MM�x�v/^�c���٪�i�W�̚}'Q�<�ҙL!�T0N�[�N�=Kp�g������|	I¼=���> �Jd�$&��O���ށ5��^��q������ݶjn߫���1�&��Z�^g&~sO�m���.�L�ա�&����@j��-z�
3�dB��5����w���ɡ~���}D��b��S`G������4D�0ï�xXlwzwZXf�2`f�X-뻨1�,x��RhYG��k=����6�Ԧ����崻V�mf�#��z��:�N���t�-]���-8&�14�]t(b��!�%��qJ�4���%\��CB)�e�OP���;_g�d�R0����t��g�g���n$(� ��'���t���>V$���}���<�l~��9�g�g�Y0��kpo���qf�o��_3��dTl��y����i�1L\
�z=�p?�dڃ�Z�$�rI�9�0��b��!'�	7�E���4r���,Gp��R�J�ȳ��<H�I�v��ո����	Z0��,�@ ����I)ZR�&�Yv̌c��3�^9��s1+���&�k�R�/Z��X#�u�[���W#�>dUx{��C�*�S�A'#�W�g��"bny�I�BG<}=a��u	��&����-�5�=����"���D���MP������F�"�R�|��m��e7
�)�3��s��QNq�{C%�{W2��hΌ���V�	p�H�����Sv*��*뗫͉�E�K�9B�9����1�H�ń��޺��T��
�~��ȯZ���n� >�R�(��� ����+ɐc0MVB�S 6�1��_v���Ek�z�����Н��A�4�����:�k�(?�Fmi�Y4!A�G����&�mlG���k���ZK�YF���x��L��0���w5{�<���+�D	75J�N6)-Xy�����+p�-̘14$%K[ԫV���4ӈ����B yv��ʽ���=�I��}�Y�������#��%	���*qWٟ
D�+���6{^�7�/ �Y+�����%����O�2oX�����b�����$Y��z+iƨm]�y��r�;�� �E�=7��[5D�Z>���Vģ,���G��EM�b�0a��]�ˤ�~�[N$��u�[�(�Z���X<p�P(,0��R�8Rq��%_ �*�aeP�Te1��&2�
��	���c<�q��g_��/W�s���8+?�I"���t)�u�s!B\�\�m��֒�³�Ǡ�Lք,W��Etjg�������CG�Ζ�M:��m�`,�d�n6qZ8q��4}C% ~�N�_���3v�=�����D+��Ah�	�Y���B&�a6��Ѿ��?E�뻮��q�#> 	]�����ޱ��ZΜ�u��/z�=�;N���UNZX� ,��d-�E����WX������LL��d�w�n�g �k4T�tW*��ONl�g����]���nBSF:8o��]�^�!0e�K��u�+O�O(&�:~n��i���n�:���kvH�QL)eCw��f�\�Pιn� `�6�nx!<uAh�=��.�Q$��2�ˢ2�/�x��{��J��z�Z�����A�=%�Z��?*M�����Z0k���Sw���ӓ)ڟ�s��Mn}1f��U�2*�63�O��X4WV"�C���5���Z�*�Xۭ���۟+�^,�������>A��x�?8�X\�"��)����&*��K����3�h��,��+kP_c�V��P���ѠY��������'m�}�x�ʄ�x��hO5O/
��h14a�9QO��.����5<XO��v�Q1:�o&8�_�W��J�}$s}�6g�c�X֡�@D���f�|�Ӊ~����]������l����S�:J�.�[j�<,�����b�yyc 7m�-��;"���vc���+��<�#�~g;v�{X���C�{�|S|�J�-l ��9_m\wj�`!&���B'Cۻ�q<qSK �e�O�,q�#������y
V0��7�$���q�t�A�ꏧ��OyqX�Q�G�k ��Z5�A�ST����pA�EKo'�������@\��AbKa!I�0b��v�ǭ��C}K�!-�_�ߘ����ej�9g'� �aVUHrZlϪ���RL�q���"�Q�͑�xq��Z��zDVv�|�Wu�E��&:TM�b9'lI0`ħ)sR��`�!�x�-0�j��}�g�m߼�È�����[��
�,��)�XYI��Yhf3�,��9��;ίC%��W�lV�Uh��c�ל���Ht�%,s���ؽ�e�4�V�PC�6_&|����R�us3<�����d��|vFL��Y,P�<)�.'p��u��F��=0/}vi�V�]2�3�~t�1ң�K��\b'k{�� ^[b�t� ��O��_�+f��������2��L���H3�,`�B� t*�2�'K�/+bIiE��/��'��:���R��! �kُV����N�7�
�NRУ���{hy�fؚ�f�{c�����	6]�c/yW�����ݧ��&�Ջ��
	p+R7ʛ6�����$m2g�H�I=���s����\�sIY͗u��k�'�΍��J�XolM9Pm����j����G����b펷zP�Q:�j��g�pݬ��[� ��R�T���7<���O5�G!�p����rgT;�P����=�4Hj WM�,� ��,%7�� %�|�Ӹˇ�j>U�8e�5����&�:��t�h
0	�����H�?b��e+V&�73j�Pc���<LI7ԕ'�NC����ƍѫ�\�G���!�\�l�:�M�i��e�!
��o�E�נ���l��"+d|�S�.���V�D����6�xG����?X��j-���յ��XA�Ԁú�b�}�=D("B��#�9O�$E�9��^Kofā���M���Tc_bɉ��+���|��h�Az���He�(��<'�Rj�U�p�PWh� ���!֢iٰ&��U8Z�/��Z)ꝥ��U�|/�ELqt�X��*\ (����B��V�J�'P3�-�uWPќ�Wʵ�]sW�=���4z�~�6F�t�]�ƽ����%6K��}�wwK�ąt{5��Z?)t�`�#r�n�x��Lh?�)��1�`r�XR]@���;��*���q�2�i�P�8�Bi�|B7�'5e�svY��ph�p��BÃ��iS�nL��P:���D:7���<0W��/[��7�	�����^�L�#�D��_�5 o|�K^-�k�P��l�x�ݶ��!\.�x�]���ܸ��͉˺��SO/�X��?���{��%�C��_��J0JV�b`qu~ڶR��\��������x9��PAB�1LQ,B0��J�lq��T1�7_���������t&{��dU��L��d4��k��u��g}�\F0��.SM���s�\+��$M=0aA:<}*"���裴���,=�ƌ
(�L�J�b�zW41aI���>���4�s��6i{c��(F�{�>�L��P�ӭj:E�X�چ�L��*6i�Q�}@�>9[��F���/��	T�"�$ۡ�:p�c����jTb\�o�&�z����p[**Xu��K3䓰�3�^�:[]	~�{� �fB�h1$,���������Q��~"�v$A1Ö������c˼i�!�hf(
ؐ���+�n*��B�u@�{̴&�%�pE'ͥ����EXG�b�&ү��0�_^�C�z]�F?{i�h.������Z��Mq\��0��U�����YN�����n=B4�S��#��q�[�p=�/�X����X��&k!G��"������ �p��ݪj�*?�Lv��`	4�tL�Z�uN��,e�VR"7�{�d���"����=�Ah1Ԟ��Q��I����s���]���ݫ�p=L��x�'��L)X�d�~��)����{�"t�i��S��-���Owq�z2��}
v�3�e�d�n2��=����Ŝ֖���d�p�S���洘]=���䇑xQ���C_} �w*Gd����{���:zH��r��A���(?�^�%�n��~ �l��k�}{�b�k�jk��ڪ*��p���и�X���4B��q8�&�uAx�K��~R�YH���1��D�P���4�|���#ն^�"�ܑ����F����ci�B���2-�T[�����O���V��w������v�Q=֢���(#� W�g��ʵ�W��)c.d4�4�_y��%۽�(Z"���i3$���.ߜk! ����lw$��"w>����Xy�7q�5 �s-��+�B8�N���Qz���Ւ�.�E�I�F�p=���w*)��)�N�YM. b�����U�Ia�S|��Ĥԩ��Y�Q3.e�iP�DC�.�vKKw��D�&�$�N���`�i�!�<�)�#���D�@�z`-y�w���F*Z�.�¢�݀�(Y1�@;4�A�5�b���{�}9d��Nw���UK���X�X�#�`����+d�̕�'���O������[UC��Y��� ���@=�Ro�7k&7��6_U��-#�K\��K�v֫�=sI���}Z�/�}R��\���&�)�'м{�+�
q1���ޕ?}/w�5-��ĝx#l��#����D�>j��խl�Ce$w���ǌіσ� ɛ��6���Y6}�UEЋ+#C��ײi��Y�b����@�S���<����3�+u���ԂB��QD�1�7M2���{�E���C<�¨dQ�m8ַmEo	�&�qՕ�8f���0��n�J@2��GDG�7y�b�\o��M����^D�~<�[����6�8�3�Ȧ+R���h%�{����e�(J-1ڱ)����/�{�ߘ���vwɉ���G$tV
���'k �!ĲȤ@���!aJ�%�Q'�:��9����A��3:~!����/�1�%Uj�
t�����o����;	�����|����(q6C�xM��@�:��C!��қVb1����XSEaWgs��WzdŦ���}�����ͪ�/$���>�4������k�=`������&=�Z���2�K��N�>�dJc��``�~s7X�'L�-d��Y���_�U�qһ�7X���o��o5�q���k�99��|��K��Cb�M~б��ZL׾w���5r�#�zq�Z\V	vѥ�W��6���{oY����E#����.iW���gs�C����N�_�_��.�7>]�LWS��9�Gc��;�SrΨ�Z��C&!�l��L)<E�凹_tl��#.z�e����ӄ�\���Fq�n\���|WpF}������6xo��T�_�7�� �?�b�kBzRy��^I��ڭ8��nm��ٻ�����.�ꢁ4����\�=��򈻉�	��ݶ�a��	7�+���� �;�̨�ZjR�Q����*��y���lDC�tV����*�@~vz�QdX�XXY� �S*nԅ]�zA�bl�����1{tI[�I]��y����ί��a�Є�s�����Vp��8A�<���/+��f9�!10��m�	+����^�<�e�FφMK��̓�8�^Df��@�m�xk46�V<��LL��x̊��yVD6a?#?JYG��!��Q;��r-�G��W.��v� ����K��S$#�撺�~|~�b	/�0����L�lm�%���U��Ť�����1j�x��W�ŰcK���.���,<vX1�eW1笜0���݌�j+�gO�*h��6d>k�_��#�L}e�]H<��/��v��/����lF���~E�qIl���i~	zl�'��ٵv4������E�y��ǲF{x���7{����[/N�;�b����kf񯦴c]�f42�E:�i
Լ���q�1�zύ��>5��#�J����5K�>Xٸt�a�aaJ�f�΢��pI���5���q��/~kw��p���p���;E�6�L���f���6!���±�qf7`U���/A�@}��&�cS�cQ%Y���V�϶���L�����W�#;�x�C��%k�g �����Y�F%���;�Hoq��0;�}��O��,N��|��P?�
���H#U-�ĭ+����*�K�M�ȝ�W^~A�j�L�D"�s.��F&Tc_!��c&��ߨL��F�#O�b��g�tsZ��hui�)���{-��j�8V�:I��-�Δ<	�%�#O�7F1�	Y�5ぞ	z״�Zl[�Y���UǸ|�	�v�$$F#c�$[�E�Ȅ�<����^*#ǼY���$8�o^�#�۸	u�>��#CN��oTb��U?PQ/��wxj"�\9�*U�
jCu0y�;>��P�n��)K�b���=�Cr˳�C�ˑ�����^ޯ�o$�9V[i��Fm��}����v�}t!u��6xN�����ml�ɭ�����w�x~j��^�
k�ó]c��ߑ
�4I�GGfY:YX������ӄqy���f��� ��TP?�U`����}' ���*܊�jYL������)����-��W�r��;��%Y�ge+;�e���{�D�����v�v��,�������޹���@8F�n���a�����&7��9Ty�5�ZZ�\�ǩ���6�Z�C�,��pk�Nd���7�k�+�Yϡ���q�v5�&�A�u�K��Zۣ�ߚ�g:E����y؍\"�]�^ ����TW�(��ǵRVj���I��ڰ�ܐ+�|om��/)'e?T��[ё��噔DI�?�&�̄@���^'�4�@�<�E$�)��6ڐ�9���&*Dԫ��W�1�Dt��H��=3��Zg�tC�8d!p2U�pp��
;U̚�]��8-��j'��ߤ�����8ʳ�����NC�;:�����ɬ`t�nIr��2�uP��w�O����-G�\�~�M֛�-A3�VPb�w��xg�!8�nn�Vi_f�9�}-��PSd�ル
gFN=i�q��1߇�,#�|>�$h�D2w�?�������f�<�M�M"���i������Qn &�e�ZY7�es�q�lFY+��7]������b��]��0�����8'�+>�����q��z����0:�����!�'v�r���`�Uľ�7L~�4�^3Ҡ"@�$ap>p�Й�i��D��QbfAۃi��I�l�kL,:�˄#��!��h�4{7.��:!��p��M��Z9�q�G�["<� �-@8�����Р�mӜF5���Jh�Ci�����gr�00=�L�8�NeTX�mګe�
9& �+t�L) �0�ƀOM�@�f�Ҍ���v��,3�+���(��y�O�q�{�u���(hKbϲqK 5�ⴾ���%s}�&M�s�Iq8� x��ãB�*����N^q�t	��Ԇ�ĥH�t�� �u(Ӊ�����5꛽�.V��X8�b'�t���.R	eĥ��]�
�,�?!R�I�>��W��L�ϒ����lt��J�lЊy�(̔���m�� _7�������*y0]`�c��׾_{�y�̜�F��b�@��5��Jm�e�:��KKt��^���+�|kaU��S���vz���A��5Wv:��r�*Q��������	7\'I����4���>��՘��h7 PQ.z�I��O}�۹G�ԥI�z*BO1�E=��1 �n�;�~�n����{X��u��،�ŉ�(nn��Q�x��=U4�q���n���l��h �[�/������m���󙗜��]K^�RO_E�1e�^j�!.��}�OL�W6�M��k7L��]P[���v�i����D�3��!_fٰ�F�H�ᠣOי�7/��;��N�j��3ڶ��n���Y�N������클٣�]������'����+'���A�����2�+N~[D,/k�(�P'�(?{зjY5:Bё�@c��5�{Ѥ\Z�KP�{R���9�at���r��ވ��6)w:����0_V3	�
�Y'i�Y�Љ��a�h*g��h>�	c���d$c��8�ͯRv�U����/ԦQ�񯛗�Q�0�a��mP�����@��rp���Dr����o<C�
����s��t�.򽉽���)�%j/��PM��,�$%�A��Q��@�6?�o��h�k"�9�{l��L2�=}	�(
3���y;�Bi��P�V<���r�z	�DhS��<������MEI�Pk�n�#��~�5^�%��ɝrn�:b��M���b��F;x�Su�3��n��6�lاm}����A���_jF]�,_���h\mEv�Ǹ���D?7G7�ކU����c��m���$��!|PiS�<;���)�W�=�ș�%�*���k-���v��	��Fh�
cA��^����&��`˞fg.d��*�x.	,<�c*,��dm�P�H���ܡ	�-B�{�&BY ���cP�5G��s�����e�$�Z����?5�f������9�<��@��I��<��M\c�YI��a!oer��׭���F�䟸�Z�?�1���x�`V�YĖG"�y��Kf��;;��!x�k�%����zo�02�^�iJ@r�j��#	�dj,��D5��؄�^�:��{�X)��!������H��O�:���M�H���0�ה�\�/�HTD��� �A��G� 署�Lh��p���v�Z�� GJ�3�EZL\S�sٟ�J�)}~y9������qgN��\K2�M[��]��.�N|^C����r��4����v~An�J@!�QrC�y�J��i>��-�Lku:u�� |��H�-�Po@$��ҝ)I�k�<|��
8;�:B������K�mE|�oV|�/8{���mb��L��(x~�������5��oo�I��o�s;UF�r(�꾈���a
4h!U�PQ�L;��Dm�DK1.��"i�R[�1�_��,!��tu�&�>4���Z��bgZ�@��KNaJ�@��)]֢G58��<�BG`Ჹ�����y'�����������3�^j)�q}�'�,�jK'xF����p<ܥ�f��uS�4��^>�a����"ˣu��Z֔�>�0���@^���ؕm�2p���6J�:B'��0��;CwF8��S�����߉����ݲ���x`/��mSPB��O��(D�XM�lď@�ج�Gx���%"�U5#��s2h� �����]�Ė���":���-r�{4A:���a�$k[�ш85K�k�[�	�&���%�$�1�,�>9�L�w���{V�g��yMfD�㣉A��N���b�4z,=��|C<�s�Șfku���gJ���6и��h8-�Ä@�7YR����+�f�jӫ��u�5����!��6W��-����h+
!��%L%�ľY�n��Wm��.�qF͊'�5�?g��BǑ��#�d���h3ezb�U"�~E�N�O�ݩL���Ѷ.�>z`]�}YW�Q��	{��y39h���Vj$��ijg�n������ m(Eg����ߡ��)0�|_H(ღ����<�ua
i����3u��XڥL�ғon}=)��w�P��4��^R�N���*Q�+='I&a��\�P��b�E�%�	+�����Jl��������ؠ��k���	n"�M6���vA�7i$�Iu� �\�c�S��Mr5,/ʀ�Z,��\�Ȟ�9���U${-�`0�ٓ98�+h{�nT�hy�S�N��������N�ơi����]��㶬k�<w*�5|�ܹ[��?��(�{�>�@���vR�����!�:zJ��y6�J�Y���F���� /kU2.���`�sLs}ՠ+e16��vB�{)��d�-ń�(�$Vf����1W���Ƭj�g(Vwǂ�F6!\�u���#pA��wp�:b;
��o�;zz�D��dSP�"�m�猍����n�H�'��b�qv��ݦIW�C��W�f�m���ϖ��X��#赹^
���~�rdd c�P숟�=I�h�:�@���r0@�Z��� P�"y �qM�%-�F�?�����-5J��WB���F���E�χd<�pY&����ֆd��O1H��I9WȀ �6��8[�l���}�y|�ဵJP.nKP��c&�Y^pk�5c��N��3[�'�܃�ޔ��ύbo���4�b[�r� ������K+�P]gA�7�Y�$+@!Lb�@a
���˂���(��ci�C��%>�9l���f��n�s�2{���-;_�xI[o� ���fV�;C�h$2�l�.��4�Q�K����(����j6�R?�m�Ya���qc�[�m�<��sQ�È�"�?�U�ak�L��ޥ�;�Fy�"�|�oMߐ>�7Y�	���7�1W%&�"Ml��x���9cQ� Q��@��ֈ���엗 |s�5}[��x��2}�����<wL�pTy�M~{�cr^r�� �_O�=Ri�5$�;/��μB���t�l����G=NPJ��w�{�e}#J��S�C�qL���^2W*n��ht���ڏ/2>��UMԞ;�҆�wr��z�� ~�0�:��}�w`c�O&��9r��� �~�<t�x�<VRD13�B����_�UOtTS�������^�a�5'z�Z(��\Z��\ٳ#������IY��扸1�{�C�a~ö칪v>��"9�5P��7$�����i(�X�.�H4�z3���Ęؗ:i'�}kC.�����I�+�6tE$ ���J��2gb}zw`���A8L�'5cw�V��6��-g`������d�Гs�L��J��N���.�`�B��ͣ6m 1�5S�>���Z����M���B_@1�	�\(���f���.�a2��\^�ޔ��e�xK�����&>���8�Z�e�P�f�Cě��]E|�bۀm�n���ĉ��C�Z�it���3�\!�%�kHIz�"�&rH68N��d���g�����Цċ��^P��MZ{&7���<�ć�[��G�-�����\�ºrk��3\�+O������%^v�4n~��s�$���و��0�"��pMp�8u.FSّ�|�d$.�����}��-*wD%oVf�6��}I��Ȑ�_ 3���/-q�jˡ^��i����amU��7�g�}X#����D<�׏G��w�Wqjf��x����Lh6����[1�95�ʽ��Q���,�]���]
�f�'��L6?#�9D��+��Q��~�1�<�Yh�AC	��"8���vB���/pֈx^�y�Cz;���[�I��� �.�<S Px��x~�S�X�f��،��c���q�3jTIV���z=��lW��t"q����C�mB���r���|��f���9��^��d��`y���}��fC���9��zJN>!�[�����#CNF���h! �n���]\��䱷rq�ḙ�^�_H@W�a|�&Sc')���\�����G-�?)]���w;Y(� ���Z��}�n3�����(��$��JF�2h�9Y��y�>�W�b�j�|�*9��?����{8z/S6^ZY|�LY�f��hϙ��{�&���Ю�����<��kS�j�J8Sm���3�?�+I�\ܪJd�@�Y���Dfj"���6c���ȟm5	j��3���:�s?� �U��w���V�"�]�ӑ�a�;z�떊��e�P�"�� %4m4xxecU��^b?���3��	"K��Ȣ�Y�ꏞj�ִ`��`<Y����=�Tfũ�CY,�U������{�L������ab��H�.I�wFM��a w�n��(��ꚰu�����}:1�Kq�pǸ� �^�w�kݘ��h����o���(���O��6��|�7Y��g"�䢨DM�4�lYY|Zķ�vf��V��Y��In������Q�<�!�Z(��K_�d8#��YN��L���㘵/O�[�����ZK�;�G�SI�cp���V�b���e��Z��pq���-�:����	3*�����E7�"X�4���4���^��4����.Ӽ;#��������:���ꖠ&�oe����I+�߼������=�!��'p[d��a�Į����`dgH��hJ��{-<�.Ż�A���Q(����k���/P]�E�oU�KQk�[�F9�3�PeR[��H�^����-���ȩ~����7��q�����j����+�4�q��6:JT�B�|H��c@��
�;!W��jЄ;6����c ��R1�dh
b���u��U�D�j�~�<��=r.6(0z�͒���n����pmOh��=������2��զ��zk��(��r��4���.�w����Q�`�T�����6/�+y�)U��؂pk��;i�),���!W�:�5c$�P�ڇ%Aڙ�����r��'RA�BgN����#��B4,�9�V%nŲxR� w�K?{�M8�P�Ob��BM�0=T������o�<�:�|�ߊ'��c��u�9*X )��F�$n�S#�G�w�dJi�&'3|j�٨0�p�h���xT��`�4���=y�p�� �ݘ��b�z�G�QO�8�/�`��o�=��c)����HAK��ђ
u?a߱�8�9��h/G&�6�u.ozp;�����j
ZB;�Ƈ�8g_��~HC��81����'��z�ި����*�"�p��ޘGxE�N���tױlZ�����3V�t��ڍ'�R��/�Ky�_������CJ�<��gM����`��:�~��U���� �5@�"	�K�t�VЬ��nVQ�EE1x����]�24�NP���qj����l�,�]&�"P�d��@վ�&�1�u�����P��x��Y���e������%''���h�=P����|d�6	�h��%�+8v:;�n���ʖ��U�đ�Av�
��v͝��J�S��ox��g�X¶��U��hNE�d4M�XM׊�O~hg� }�;P���L�Q�!?S�����|`�����Qb�s��P���7~�OP�l� n9�6�#�9���,у_�^@�*p|�P�x���(�ģXN���b�9��uN� C�o�Π~L5��΃�C\5J����5��Z	2����_�`F�t�,�t�z#��h����]k6O�"ךf�"��x^�DEKB�A����)aa�����σq���[������ӭ��Z+��
��݄N���%�������x ��N}ߞg��� �/�=���jb�z��h�oo��H��P��$کAN�؄q]$9lPP,ظ��3-RrʟB+�	�i����C.f]m��zj����chu�Ly�>����+,�l���6��/ݢ�pC�L,jZ��N�m�;�:aԸ«��ǉ�W$�_�Obx!�uՍ��͗��p����mW�c��x�o,Ѯ�To*��BW�4X*5��S G�I�B����n�#C|B�/�8�<����n�XZ�W:���䗕�p��K&4?�R����M������4 ���Ra�Sm�Iخp�<��ia0��a�8>6���Nx׬Ӑr0ދ�ؿ˖�����}CbV����V8P,�|�Z�co���H=8���ǊM�R��<�zq	��2��� ̹���;�X�}o���J���}�xB���g��ql��ְ�����ꐜ��A
&FPX���A$��1�D�W�i ��ܫ��M��-�A$��S���U�d���`��B��]����>�[e��F��be�&�i�!1�2:�<A��b�ƶ%�����f���l2��sї��e���4
�X�}�X������V]�)��=�c>��8wu)���w��|��_�~�kh���[G���D���>��Y	�v��@�k���	)o��g54�ԩ
��Z��tu)KtbQ�|ޅ�a���r��tq�C���qM�A�T*�	��w��*E�3đj���x񣏥.�)C���@��`��4k�T!�>^�?S6"�?��������OW�1�B]�ъ+���ϵ^û�W�G"�C6u���e(ĴJ[d@�ņ��Y�U<�4���^�6���7?�X
7���y��zV$p�˰���m�����L��<.ݺI�{pĳ�P�G���/
o�mvZGX��w�xvD��YQ��>���J�o'�	<�3T6�����_2��pl�W��������\�C=���g@[|͐@��ܚD%�W� �\�;�q��N�|�+X�Vt)�hM	db�)g � ��v2���5���I���	�"J��vp쳵�O����{�UO��"��G�7ه>��;!
o�W:���4������ӮI������rąpo���`$�����LC�7�0`���������#E-:�lAF�tDT��j��B����u�i�
�k��(PhP5�!���(����X�SMz��r`Oy�rs�j#�Y~��N���a��
8$y2e2E1�_�׭]Sv���l�;�D	]u_�C���8G�HQ-���� 1%] ���[�FJ�y��� )�8�$���g�6�ܛ��c�zG	 �╙3=�����T��� ��<c=y�z+�9z���hL�2~.�=$�!���Vm�V�"Ud���N�a5 ���1P���a�����m|F��c�d�p��:Lc���nNd�Za��{-�[W��00�NC2w����sȗ��S���� ہk��y�����dʶ�i���H�I_�������*%&��-��8�'��:,��,L��%ht�n��V
�a��ް�"�����������6�dwJ���k�\ �y�ډ��᭟Odz�ĴE)?�yV�g��|Û6��Y�����Ğ!�s'7{<�чB�9\��Q@X}<m	f�oEG�	�3S�����!�ubOS�
;�I�!UYHN�G:k�X|
<�7��2��k�y*���J�H�����p�A,���&c���ۏ	�W�,�0M%=;&�A�{Յ�4n}{�5��`
j5
�n.�XS#�~e���ߞ���!��̏0�$$7J�-h�C��n-�r�-	�.Q,����e�� 5ޡI��I�#��a�5L rhj��zlM�߰�B��vP/I.8$*ǽ<�E\T_'�B������I��As���C�&����}������o�{��i贄�������~_�18�FQE�/�!]��o�i�Ya�g%# O�0���՝
�K�(���q�%H�U1Iml�9��`�=�,�]@d�p	��ok<8ޢ��c@��X�eV�Ꭴ������⊯u �h��0F��3F<��Q)䇆�X�%J��ݖ��S�?z���/X�C��$�����={��" ���{�A.�{��`�6bdܝf3��O�OT���a(�ݼ�T�s�i�=
�����N;"�����T�E�q�@�C�������ȃ�ŖP8(F�jɨ>�$�3�����:���c��������ՙ<�,�ɳ��Y�߆8ӯq�֩��g<eWP ��*�!���!wjd�^kT�	�T':�0���)>��)�-�Dte�H)N*��g6�������w�~v��W�̳�`pI����O��������<U�ܱћ�?�lj�~�\	˛Rx3����|�I�#&Q�I7���/��.��g��p�����Y����pw>Lo�A�b�[6��5�s�7�x%���VW,������X3��͍\�8��Q!�ԎX6[i�)#�����P˭n������񼆬�q�H:����vw���Zl2-sIu��Y~?��A���8�)���n�uvc�"qv�F���)P��>gG/:����˘���L5��*�߯RF�������  V�G�~/���ÄW��46�Ͷ��Q74V�X�n�<�1*�h)�'���Kc�"����<kI4(��?��k��N�՜����T�7�Ʊ������tc'��p��L ]r�9�y$(����!|y�������!ֿ�к�dӒC6�v!lIL<y6�
���TM�z�	G�h���}M�ؐ��y'N�J8F�)��X�٦╂���~@�;�3�ף��uߎX�2gB���=ZȌ��eDx\��WJ���Mb�� ��I�*�܁j�#(�н�d�8���6�	�Hp�3��J�m9�"��p�UL}o�^J��U��-#�[�i֩��j�E�*J�"���'�w�h�/o�	;�	����p�d"��h8�0�1���@����M'?Ԓ��,���('8/;���r7W���q��A�c͋�eC���~&��B�(�*��m��PNy�2q��f���s]%b�PʘT>�0z��1=�����O?�]��}O/F�*��1�P�H��*��3���̲E2&LA=���ٺn�b���Z�R��DQ��4�-�'���jxR�� ��&�����ȧ�C����UO���2�G(��uqz�g�_��A�h��Y���E�j:�X�jU����Prj�L���h�0eL�b��V;v��	<��4���\�I�1���w���2c���(i8��I8���Z�7 �^*�dW��;�2�2_�j��?� ��߫`���j�Y{b@�Mb���ד5'�7p.#�Mp#��`���E�bX!*ߤx鷾�-�=�=��'�7�G� ��'������X<��!e:�B(����sRt*t�r?e�k��M4,�r��U�5b?$�ˣ��$��Hc��ta���z[.���k�j+��\+���Ɔ�tKccL�|kf��?�=0+�'�zjQ�5�����F
��K�r�*��x^����S7������*;��b�Hu ͗�rff�R�jK<�w����{�Z�F�-�L��/;{����3����%�o�ux�>��m'a4<X�0�iɘ�1��}yhfl�b{x�G�_�.|8���P� ��<
9�]fz�0ʂ�-�Y�:�������|R����6QȔO��!��|�,KfeE�,`������VbƤ���F��~H���A^���4D4g���:�4hכ,�����e{�H\�U�����n�����WB�˳�,��H�cj�)�6����z�3�J7Wō���U#\b��y��+�ǅ}z�v$72�aUM%:Y(��l��W�jh�;6�H_n�d!,�_�|��<ö�뵔;`��0��I*~�nb�b����LD�V�
�h�BlG$`M��j��v���N��:�z�f���\�Z�nrU@.�S��,\<B$�o�5�u���@���,����J��7sVڕY��D�j��w/����[���X����������|K�q�aQjzB/{آ���`���݄�nq1�枿(�8��gu�\*Z����.~g���Fm|�c+R127f|%���u��8�
K��������{� ��0�pw$)��b���:�cpC��5��l���3"�Jw�7��и�Pv���8�1m����{������ΗZE%W~�����ky����HL�q�ٕdQ��Oy:�K���7WO#z�|��VIT�y�"�q7��/Xd�B-��~����0�2G� ��S�ク�#�=��XQ��l�%Hl�38��B�,�8���I� 1v��S�xb���3� :Q|Í�)�%n��ѻ����gR,m-����&�G�R48X�Deb^:��+��x`����; W�m"�iZ) �W�E]��E�g"<�ה�0��l&Ze�է\Uq�9o������թ���C�~h�������I\�`�VM��]2v��ba����|[�HM5�,C����d]��i��*}sK~�'�'��(K�Z7��<���o��S�xJ���
3|�9S`0p�Tl�/&��^|�y]H�|	�I; f��γK��<��r�=	�y��)��g����J~�������n�*�l�����y�7��֋'�,*>�ė\�"P����V��2�E����@'�����Q�V�\��Ś�[�"�����	�,AS�~MK�ɚK��������V�������!����M���`�����ԯ�a�����d�A*�|�)�i�#�����9N]S�G�;덓���4����V&~�G���p]���|����8cTTES�z������O}Q�����VVۮ1Hv�޻���������p~_��i�U��e�{.�o������[���QFn�M��UUc�K���7UT%�Il�#-<UuOL%�H��C�I��V���>����nl_�����S�V�T���Ԫ�VG�_��d6���ds���֓0��Q}������K�G�ԁ4��o~��E�}�ߖ�_I����.�+�5d[M�	.��ح���i�{G���q2.�Z&��i1���S�3�I�v)3��òs�g]Jkx�zz��uzAW
��k��G�:p��uε���K@�BUG�a��8�ǳD|P�J�D�8'Hʒ�Vˈ�h��:�3O"�`r��.��N�pNW�Vb�F��|q��b���Y���<��mq)�7J����|ԯw��IQ�����<����U--�m�z�4$G,����:�`P�%_�1�cĚxa�2=w=����@n>j�tL���oƘL,����,��_��q~(xU.r�o������I	�H�������vm�^��JM�1�C$��c0�Ҷ�;��m}���k�1N[F5ު
u#�zm��QiGz*^<�
��L� W�����K[ؘ������W?���%bd�O�,�	�.ł�J�����]Wh�cט{��K�c����=:�p���^,�Q/:s��Ҧ%����М?��%#A���xB�h�MR�p¯D�,ɛ!��G�)fpxԄSqR��D�FzHuO����׿b{��cQ��H�R����j��kF����]<Y�q�C�f�d=�&����Xn	�+e�Y��0v���x�4�
fP�K�\���tW]XB��7^i4+����Rt դ�+l��+�l�(m��g1-ڑ@�Xo�������c/?]ܰ��:�ʿ�	�`�w�s�I���.������ii���O��f��/a�+@��q�hz��0�u�X�&'�6��R�Ӧt��>,8�˯d{F@P`���� "j����干;{ƕe&�h4��W��K^�}eM���u�4I����+P�#T��~ϡs��qS#�צEI�E�Ǎd�L�6}=�Ok�Ci�5���S�|ㅻA�H!�>#��v:��v�-W� ��Bә�jq�
 �c�Ό�~;$uň�z��̓�?i�fuF���(l`x�@�u*u*�������k�K<$�k��׿^Z���jH�Xf��I���1@e_aoK�%�_�V>��9��3D�sԜ�k�	��1���a6g�n��?�?�8 "Ȍ��(�7�s܂����6i0C!�/f��syhK��p��%��]��U6���CT���և��|�c�9��bߏ4-.��?0��t���G�m�+��Ɣ��.�`\�V������s;���`��8�?��= d��~�o����4*m`ǶW�"(w�09 \5zLT�Q��'�l�`lQ?�8�#�E���vn���Ǳ$Ľ�P��o%�j�n]�:ׁ;:���M LӁ� �_�ֽd��p���ȧ�A�^��~�,�s N������F:yIV�ȗQ>��ׇ7�c\c�)_�	i��ے��ɾ�\ٗ�j,�fw���]��r^��Ffm�:o&rp�!�n�S�J�{@:e3�'�W���x�a��ʴ�e��{P��G�)}M*�,-O�Qy7U�j���D޳�ѐC��`ͨJear�
�OD��g���{��4p8ceI�=��ӻUQ,�ߠp��^��q�{ŭ�̀LF�mR`I�w�B�����=���i{�\���f����k[[��C��z�C���r	�(v��N���Z�1ܥ��}_^R�G*b�����Ċ�1�⦧��~.f*b��[l]��Uͅ���"QN�o~#���+��~�_$P�ی^=�W�����*LH�>(�ҝ1\����4�ϒ�J��E��zvL��(�'�c����0��_�yYMɍuQ�3,G(?\^e�����?��ؚ�؄Rk�:_�����+mAl��D%�^+l��j������G��n4������Y9�h�Y��b��so�A���|.L�X��v�J_�����.�����n8���0�V�y�Z�EJ�N���/�,���,}U) F�i�
ׯ�@�no�0h����fA/&�3[�����(dڀ�����嘟���>u��;������G�Mf򺊕���>�r#�ڐ���<k8�d���A��y��¡*e�8�w�h����ʨ vo����.����o����]Ek��6�Kb=J�Rފ�.LJ���LՑo����*J�Jb���>��~��}�)�Рx|b)i)�=����W����Rd@�֦�8	�o4��W�Vl�)u��n�� �I����0>IW��C����v
 }K�͒=��Pe�Ѷ!섒"���)
k-�p94Z��F.���0bmS\�Pm�ƺ��ۼ+>;Υ���<|��4ƽ��WlA�f3�$]���{_V�E]�֙a��J������=�Pvc������m�洸��U��7�ə\���+-��Y���hK��D�s|c�Tݚ�{l ~u��n	ԋ��	�F���?Y[�Ć>!�Xʆ���1�.%�����	XAtVsZs�@��2T�p@�����H��awrI:�ӓ��BoX?坯��(0A|O��k)��F�W�2�X)����ܨwQ1�~��(AWɚ�C���@���|�����j��(�@�{�A�B��j�VH��Q �Y������^�c98I<�+����
����1_��n�G�/��j�Q�[��#�]�q�2Q��~�A���
��˹�*�:��if��0qqD�5���'�:au+ro'>�A�f�z�D���k��	�@���b����K�J��Y@���Te��=0�R).���#u��eO0ϋ!@���� ���V)��d��{���n�"��pm��Lg^�c�b�Y~3j�2+�
P�ض��7������*�ӻ2��j� O��yW�]��i���ts���f��K������#������mM;w�)F����zF�d��c=��q��Q�H��C�֌� �=�X��|7���@@s�=HI��|J�
K?�>�ee���}e�Y�1F��$lrE�	ݩ�(�j�����w���u�<�z��+ֹ�iE�z/��%�������讵�^�u��v�
��9P��"5&���[ǔ|�<m�2�U�����m�N�#!�>)��d3�&���駹�P����!9��S+�c�w�C	C#)����y�$�i���g̉�ܴ)�r4��;�Q5S�����pѣ'��}��k/:��W_���^] c9<x��L<��)L�vL�?�Ѭ�!`���j~H���5��d��y�Y�0vq���'n��Kueo��|.��s!�Z��EH��B��ϓ�	gV\
 ��*p����R5H���	�ze:t��K+]���34һ�y��8O��Sw�z���j�?[SBw!CmV�%u`��h��[�e!9��[�c��P���H�Z�_ua�߁�k�j��N��a
z�!��Ӭ���p�k�8h�M��WB'�L}g+���*nX�
tl������Yf����C��ĉig��h��3��x��Y��4J,�'k��c�A{&��c��-��v�q�GY��rm�`	��=���I�-��y� Л�B 2ۿ�&��3U����!����n(�x���G�o94��  A��0���[F��4K�\���ĸHl�]/�-ta�R�J���!�ZH�ȯ$�����m~�+~�S�v-�+f�a;�Nh�u�5�*5���m�����ʥF�w�����ުTu���d����̌V�ΐ-������������+��d� ��I5���=A�9���zύ���)���N���������3��Co�F�2T�Z.ק�������K����N-��
VgVF+�@p8:W)��O_X��P�Q�/�V��hVc�D�KW����Mܵ�]��~-�����ҕ�rM.%�7l&N;�fSq���}�o�m?������D�\5��L�V�I��~����%��d�^�`��}Gs���!����k�X���}cݭ�%�Ϲ}�r���{�����hZ�u�C�f����j�"�W�#,2"��Toi��eoµ�S�c�cϞ������̶䛭�2���]���F�]�=���3.��D�e�[R�x:7ɢ�%-�Ŷ�w�{l�;�i����-݆G}��Z/Ȯ�L��4�%L�V�"�`��x
�}o-dQ<Dز��T�f����ot���1Hٸ���v��)F'p�o�eHXV,R&N��A
�ż�Km&�AD�k���i�}���기�q̨�m߿�4�D�u�In�GT@�X���5��q�^v����\��"g�F4�j ə���j�&�O�ej�Q�v�)�R��I�̥Au��y�p�99:�USD��3yA��nd����I���iH} ��~����m��B"i�rߚcrAz��/N�
�ܺ�K�0om�9���@��X\���f��]���4E��ުp�@�X�$_w�1�T퓩��H[-cb�X-e�;=B�V������[��җ��,{tH�I"$�u8�$ps�8E�LZ�\��L��$P�I]���Ff#@#���|H�~H��e�~�ɒ�`��Xf��؁FE�o��+����;��1"�0�?��]�N��[~h�a3�F Q��}�&\����v> �8��Ba���`�$g�,!�-{����uM�0�I�hd�螠'�3�$2���u�v�ݣZ`]��9�{����1�u(�o�H�f���o֥|�{����(����#��$;��6��;F�|��NDi�O���Oy[y���ٰ!����z����3o&D}c!x��~k�)�\/�ON�s��a ��&����S�r�fh��Đ�c����_2���m�Q�wm��R�&U�N�� u)"R��a����H��_Y����^�:F��=�N8FD����􌰋d3�
�