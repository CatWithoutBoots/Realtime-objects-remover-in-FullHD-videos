��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P=V��F��~����2.�r4��:�Ŭv��E�I��u3�;�"��~��}_�c�d%29��H;۽��#��DuNG�ħ��/�?��+�iZ����W7��|��x��]�*d�Wy���7�T��Ez2L��DF^��ɂ�q"d;V���ٮ�E�uFI�\T���`�@/�?�rj���Q �u��Om��׮�h#9u�ڨ#�x�0ޅ�6]����A	a�C��	�x;+@�g��'M[�bӕ�Q5/_ gД��j�rא��`͎F�Jz9Q��U.�r�p��if�H�h��5J�1�]B�ьJ� �XCUY�<��7�l�8SMh����1c����`�B���:�J��t����yt�WQ��OT:<�}^U���eX�6f�t�Ë�����[��$^�:�K���UDE��!��P�i�7<�H����r~s:�T�z\��	��Z�����{C�׹{.�\��4�ف��}D\2�wTq�?��ozc�a<ІD[M 5��(��"b%^��w�n�ᡱ����A�J�3����B���Ml�g#��� ��B�����3B�x(�����T@�B��[������Ii��S���QfX��AӇ�����Jm�8��E*Rhɖ1珞*3�㲪X`�
�n�"_/Y�I`@N�{�K�K_��A)��7�\W�u�ll2_Z���W?��i0�-������Nq��[��4P�Ϛ�r��<�<���~�����[��s�*�Οɘ�`#�'�{)!4㯷,>�o(#R��
Ϸ��/*�l�����[�U�Kc�N{���e��=E���ً��=��,d���7I���C���jo�-����W���wBEm�l��o��:e�#��"vf�{|�Ғ�$�^X�#AY.��z�e�����a	�0�07������-����t!`�[�4�D�>�o_�����6 r�c݀\��g�����w��.��Bή&�>���/S�����Ƕ�ګ�6�y�ge�T#� nK�'N<�� ����?VV:Exo��tqf)UYz�k���2�+W�V :v�vrR�����0=��n�O�q��.�� d	�I4�~p�\D�nB��50�,��x:FD܏�s�dw�Z�4+J]�n��4��EI>0F]���� N��fw]�I)*�3��#�AL�B���e�it_0�Y��pV�4/Mh�	xd)̲�A����@<����d�c1�a���0���Z*��z}a��p�R�x��"�p�R}�Jd�O��^V�kDǒ���ʗuKǒ�ȹ��!h�W��5#�H
�fD��j#]8�50�.��
r�Y#:�7��մkC��/A�J�^�8+]���&Ǐ��!a`� N=����B��mqO���;�㪬����d�ڛC+��{�&3�Ho'�@(�=M�9#;�e��B�Pj)N<��A�@���r�8����b�z:��M�,������8��lo���m�i�L~�K~��Sd�z�S���,�-�j�� �`��Wr����{P0Zj��v�u��p��;�_}:R�, t�F��qn�u�֎U(�M�*(����bE�_ ���������|A?fP�M�!d���<��84q@�4�C^e�iM'�dgU!}�k�L���{K�k�I�<l�v�wM���{�%&�@�Ci=�ɸ�7�Rn5��f��{X��Hg2�6+�#UB�,Qp�vP��E���^j�l0o j�l(�RsE�yE��_P�!���K��bAv���
fи`�@��]��M	���}��bX�����;��ak�cX�&�vI%w���v@�{'-��mf��)rR�2R��6�!�*{Nr�,��^2's��χnT���ӵ�,��}���NU� Ļ��ϐ��G��|maf�Ba����\��y��I�?z:�ØI�ێXUO�:F���
�oBNNgu��g�ƆZ"`v"�R}�+�j�I��S��8��3�ba*,�)��aO	��MU痘�:~Yj�}&I��y@ac�>xQ�G�����8D@�b&�+��=u4���ŀH�b��ʚ�[~���ʶ=]J(�O\�s�kF���җ�1�4��F�V��\3ĵ3��e��M,�Y��LSo.9d	."i�7?�IF͖��ؿbp�G���2���/�L�S"�q[��}��t�|��ʀY-i�>j�D# ɸKu��Nf=Q� nl����$�Hm+���@��È�e?m4�k�@�l��7X/d�X&�V�g�݅�.pd��\@�
��}�屭Y�.J�t,�m6q��5Hg+f�V�rph��d�p��m���m�t�2�'�D23I��?�5Aİy�X���ȊN8m�����d�ڕ�DE]hԡO#�myo�_�m�_�����r�������Vs�ٚ�P�q���u��_�(���e8f�����i��S�55l�9'������'��4������TF*�t���bT�[�V@Ec�.�#��"ѣx�F��jk<�,e�����O�s��fz�E��Z��E�����I\�p�xj
:�S�
�}��=^1�� ��&��{{4 ��!+)�9��.b{��u)G=W����m�9�F'���*A�J&��
5&؆�Z����%��>�Fõ�L�ۤn_�+D@�Ih�@�I��%��#�59Ml�����{?� "/N&)\օ/i���om�%}��(�=a�K�p�3����8<o�(��4!�9Ҍ���#Yr;H=TP'/rwx�H�Vw�� F
��ГF V�EnV˺bRc��l��l����<y�V�onx9]n�6t�;`���	/�KzM��η�ra������	0��UI�x�da��ۅ<��K���ƻ�w�XM�
�o%I���!����g�)�ɎP��
s�X��)e���nYR����8������2|���������۝���,�G���	��k���B��Sy�U�#-I��3�������<��
��]0 �^	y&8����g�����TE�~:��- ��K�.�v��h���oZ�f�G�j��cO3&����sx��"�����$���wַ��o�w��´�g��~�(ZN�Bs����@|�W�%jbw�&Q(�y4��?�|��!��H�Im
c��h��u�"�$�E�PG7����r��E����i�#�Xqu�"��N�`�@��\(��v��s�3�}2��˫���L9��KUH�]���RkP�$�ܶ���31��M[�R�F�Ņ��l<'�2�h��{�� T��Z�a$|ڮ��0*	�N�c]�B�q�1k���	y2��� 
0�Y�Jd�S�G"�5�QNsڑ��r*�{d8�4.��|��_��$�'G��A�B��H�^7@=��	���|��D�J�W����iL���o��c��������(���u��id�!��ā�6ئ�[��S��bl���S1MT�{>��NC���GtK�g/���.������w��b����{�������QC����x-��hﴠ�0�)�z���9���qy(e��\Ư��v�޳^����� �n�e�q�I�{�DE��j� h�l�K������s��Z��[P��u�%WvD�]7�!(X����)ۺ_#F�,Q!*'����P*����n'wZ�$;I�1�Px+Q3p�'eN$���Y��xY�GLN0�7"��Fj��	�����'� �sG(Y'5����"k63j�>�r�A�KdY���c��#8l���']d�`;���Y�j��8G���r,��3<���O{&1��	Jx�DO7�+���E���l����D����V�d�����N0d��Q�Oƻ����N�z���[%� -WLح0�&���t��P���0j7Q��֌�Z���\�|
����_]sә�Y�L����T5� Ȱ�Q$�-�/�ܝ6��\f��(�-��Q#�O���Ь��YO�O�3�x�� ��W����p�#6]O
�*H�N�a�� �+��˸��mٴn���	�h�pz����t���cc�_+��À�T�� Q*q�qJC�I/���ݡ�z-���]�WUh�_�XQrh"-�@���)�yQ��-�s��?]ga��^��dP
d|�1�n�63��λ.R@�M�
��.fX�P?c�S��wt?��2p!�!�Ft��gZ������v`��{�Ylq���
�%D���{�*�Vd̨���/��8#��*������q|<���3׭����[V
��iϴįΙ�x"�<��T0�}o��5Ku�A��Y����󩪁r��M.�:�G�)	e�;C�nSJv}XU�����gWM}[��$$�wa�V��`�I	ӱk��堌φ{\�(���?U3�� k�Ȁaa��.����@�y(R#�K�~3vG�$TZM����||{ã� ����'�-�8��=���>Lܰ��x��ۭ�{���|v��CL_zJ$ ����^��!_ǥ����g��A��7w�/���ጨD���TN�!Gː�W{��##����YCD���o�'��=5?�I&G[Ek]X��,�1iޔ��!�ү��#���Ol�V��_���tl�����u{�����[C0��<*g�<�_+A�H�6uH��^Y4���E���c�_�rE��/���ya��"��9�h `#�i�͆!�p�����%��
����($�R9�EJ����A��7��pF�'\&sGϺ�ͫ�wH��X)� �z�����'=F\�gm_
�P��%��y���~�/���1�6����-�7F�J}g�F[�Ue��/�Z�3W�9ݳJ7�0��vÈ�mfwd��"w�&#�'��Q��V�JP��7"���a/F
N��r�-xޞ�^Gg'C��fs�L��of?ϐ;����6����R��0I�!�^\�� ?�T����2Y�®���C0��Y�^��I�נ�BB=p����3"@8�v��T���?��B���Ҟ�bO�@�Ql1ѽ��6宭yZg=2��T���I%��W��K�@�ռ��#�>s�9'o�	�#�4��Szwm[���"�墾*Jt�\c��TY�E��p>yڤ�U�%�٦�i
̪G>�����Y�A�w݇[�dS]�p|����ºMI�Cm�d���&��*J��mg��;2}0;�"~��� ��eY(�{���:s/�c�f��������|�|���������Q��wY���vj8�$��<��J��.�����"�S�?�l���j���j��}><$F���b�$�,�vX�$�����0�Y��{4����Ce���k=�&��'���"Ӵ�3v �zԿ+��!�iE2���l��hO�p��e�R�<�Â������來�	�	�U�7��2ZQ�AE��[;���k��V'�*e��G��b��s�B5lY#��l4�o���P�[�<�����@*��i��a[�s)x�uV�L�H,���g�ʉ��SVy�n�Cd�Z�eA,��$Uz��	���)�Љ�����X{z3��.Ui��,��ӓ@�sY5D��H�@h��H�2�S��7�&]D#���Qzv�$;�f�I%ϊhub���qE�~(�}c~U�H1_o6��7NT48��Oea1��#X)[O�?ŕH܈֙���0V��b����
"��XQI�`�uS���_��-68ڼ�&>�`�9����L�^�fŘ<��u��1��#À=�\�T�ĠZ�}�u)J�1��B�ᣌ���3v�?�-)��#�i�q��bq50���M����'�gݮ��e^;��	�?u}Ot�~����|�Y�l���,G���뜪[�+�:ܓ��L}�h�*5�ǉ"�9�� ���Eɤ�:��`Di�e�:��}���3�3��*
"-�]�;Q)��B��rUb5bJ���m~a�*��|�\T/�=ZuQ�����W���9����d��\�)Z��-��˴˨~�9H��F{78�I�hp�˗�ؕ�����L�]Y��?U��