��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&r�F���oh���[ynnf���6_�� !��-��!%�8Q���"�I�}I��F��ft_C]~�	�=j��)L����F��.�A��z�}藦�|P�eU49z*���z�^m�؝����5kq��>\��#SA����:bUV7�օ�>�>�	��������� җ�1�A!zW&B����Ld�� +����y�:�
	�<=k�_�9D��;��dlⲳ����}K���|u�����R8�Ȟ�����#]Ꙏ��?o\I�X���:�M��_]�n�:y��xQ�����@"(� ��.�V���0�K��|V��g�<����44I� � ͐���啚W$�~��-i�<�(ytoT���L��@`㋻�_������>�ߙZ.��f��2`���ʋ�0��(�\]4x�.k����
7�z�$��8y ����s&���ʩS�'�K�@&>¦x�
\����A��[)5��ڗ�

ЭQ��D�c�ܽۇࡠip洼Czk��x��MJ��U�(#�]��>���g��d�)��`-�z3�RY����Ღ����*�	E��u�⢬��R���.'��y��!��U�$��ɼ�1\��%�=>쑖u��J_k��`9w�oէ�%�%A]@�ӛV(d{��J�X7A|�R~��z߅���ʝ�Z�6�9���bД�?����V�%k��mWS���v��M�����K�o�r�F�|1J��������1rn�� �׌�A(	�Y��x�w��Fծ��*�B�N	NSo���z!��px�mz ,�H_��%=��aFno,�f�Аi��1��/Ѫ8���JW �O� �Nj����X�)�}�M�F4pw��F���u ���zE@Q��xoM+T�yY��B~���5^��+����f.~ڙ0	��%@�m��hSֈj	��ӻY�3�ò{��:�c�T��N��8�</0V������J�T��/��v� `�`!�bb�ݨm�S�j��ik*�6O|�՛���|7�c��.���#蠫e0�w��s���&����q�FL����T�| ��X��zs#p��T�b��Rv��!�/�5���7�`�,\��H��󐫨<�v�+��� 8gQ����6z��J�S�����oyD���:ep��l�Lܥ	���Y٫�_Ђh30z��c52��e2l�&�4;T��PxГsP>����ί-ce~$��_Zn�5��F~��Ү��U�F��\;O)�l���q�Te�.�N*f���w���F�!P�&�dJRu�`}����B4V�<s�+��?�g�m'�!O8��0�整 $ю� ��#L/�����/vwN�4dQ?Xm��2�B�*��[,z�e��7�����r�ض ��+���S�NV]}2�Y�S
����6\[n�K衫�����V��f,_1f,�.[����D�Ø���8��-Ū��]u��L�_̞�n1�-6��^e&#J��%�2�-��Չ�T�h/WK��_'�
������|��x�-��w��v��監�?Jg���?�'s�P��r�Nl���Zo_�h��%�-��~���`�������L*�ʹ:Y�D|?ђ8s�v1H��\C�1���@���7�	`3��OR9du.�`Km�>�sln�[5w�U�z��9�����}��2Y�2C�"�֕�?�=δ� �1!���\�rY�7�Y���{��HW�@?w�Xn�7���:RN�yϋ2U`ፊ������-�cG�'W{ �%f�"u��Fwn��pN�Ɖ����:1�\Gm��]^�Q�إ>�@��W  �����;����C�X���Fw �Y=�rÕ3���������c}N�
ȣ��~�s���ms�V(�_�3*���I8���A���U`��A���T�
�po_����� pu2��N,�y��`��r��Tc{�T�\��Rԡ�sp��v�Ab4�)�k��C�ݦ`�C}�ub�g�|�g��y���Ӈ1����C�\O�6D�+s�p�LR�! ��5�ZK5�}���$������c;��R���'�,��w��*�xx}å�ʋsDzB��.9�֪n�>�p#�U�AÝ��~�8��x7|ȥ 
e�8	U�p�ӨC�8�^P�8��i�ؒr��-�*5IlH�kmeq���N�p�K�|"�S5E�7� 6\���ة��&g/X'��f����a��O�`���X_;F�����`!'� ]� "Z��B��z�+�=��Iú��.�S�qe��zm2K 3�&�9zr�<���8��ViMV��h@�vO����%�c"�}z�V�KkA{{Xn� ģ�G�Q�g�C�.a�Z�(z�D�ɰY�
�)�w�C����1��[����R��,k �4�ha��W��L+>�~j@ Ad�:lU2� ��$�7������~���S�&�:�4K�c�z��@��is:`��;����@C�����0��t�;f9z�dH�p՟��0��J',�k}�PY@���T�=�'t�.q�j49�U������z?'2]���1��'Y�t�:�Ozة>b>V�$8m_�r���6���|�e�����e}^� [���%9��o\̝���y!�V��4�Q�.k.8|}z�'�LP� ��
K�U�gP}t	'(`���"S�2�(>b3�ǁ\�3�{l�( � 7��Îi�[��9�D8֦��E�qdw�]Q>��9^��!̺�6H&J���4OM'
���o=���>�@�+Az����ڨXD�ck�B�00R�[��B�:�JL��W[�o������G�K���󷜗]#FS]�W�����D��� �57��u�E�N��[��k�:�R�[-��Y���I8P��6?}���'��vK�k}�OOv��'�.��Ǵ�6߫Iӌx�
��r�%AW7B��ʥ�A"d�O�j����n8:7��w�3�/1��w�k�/f�<����-(Gs��ܐ����/�N�]ܭ�W�%BuO����s/x7w���(y;�i�ٝHg��Ô��!����;^�ꦎ|�m�=e9�mGT�V���O����&1ytؐ��o�d�~\E37SV�Sv$<R䛫Z�,m�eY���\�����<�Z�
�`%�.A�,���o���5����b!#-,�S�q��n������2��*���7�[��[�?�[�PaWN�����$cn��g�p����<���W�Q��j{�{Xg6*�dt�j���Lf54�#ɽBLC����7J-�:#���
z�Yu�[��:ğ��
G�-�~~k�>	@ʦ����&>Z�M�⡷�g��W�Ė�W�Մ
b�irҶhwO��<pD0p����k}��D8Q�	|�uy} I�8B�f���X�>�82�t���L1x�Ǥ-{&;6���0D.$��<�ʎ5�b4��1�%5��9���RW����2^�S0YJ�4�S�&\��t�vp��ΩX*{�^��+��Ʋ��z�J�N�j/��}�������<8���-��'�M@f�2��CIk�@㒻�}^�N�d�#:2?W��%�rg��-�;Idwq����nVsk���:XE�E���h[%?�KEh ���X��b��(�٠tPJ.�+�[�d��ʁz�T�pa̢���kgDr����]
lyW����ƀ����o��AˬZNn$r;G���J������,��G�����>¿H��p�x�������.����&����R��יm���r�a��B(�ENT}��dM�:��:�P�'�C��Ut�c�%=�c���?z0�4Yn���c<���I$r4u�U5hЋ�{6ۑ�h�c�<�W���Ǽ�!'L@�1:��I�j�4���`|l��[��v� �������O�k�B�k�2��
�ԪŠ+�;����c���*�22&�Ԋ �K��4��H�uZ�\(��kj�wB����k+�U���d;M�������X|Ѱ��SM'ȏELs��ake�Ol}\ãY��"���9����w#��w�M�5
�swH��o*����$��&�z�3��t�ӊ�|JZ!���l��ifY��nϋ��U,�W�(����[�u���7�"�����O �j,�/��c�]���,�e���� QK�5o�9�����	Q�P_�U�j�#�qy���/�����:�S1_�j#x���@ L��h(�����x��U�g�=&�P��c��
�a����x)������4�ƸE����=��"ɬ���Bǎ}�MGޕ}5�:z�9A���Y���=�qqxްmM0"a B@��t"H����1�v c��|��aj>g�3Hl���9!��b�K"T��J�G��(��܅�3"�����۽�3��a��f+1�jb@}�!1�3�;�T[����]�����8V�3^���c�ԗ%�(�	�w��.��'�$h<�CB<l��j
��3�.�F>�6ސd�؊>{-Z�9s�f}�{DP����H���"#�?\#�����ne��R�P
����zV���f^h�e{�͹��/\d���8�.��ٿ8���G��+)tP���7�k%�B�S�є/[[Xs�\��>o؀f3�����t�c��&$��w�16�hE�U�%��5�����}u�@%�-X��/'�![�Gcp,��w
�4�Z'����E�i�������,��S���c~Bf9(@s�/��bY�E����l`������GIZ��?�E�}�) ?���?F�qOk%�v�[o0���G�?,��N�k�!��3Gv32T�TQ�H��i�UW�|p+��R�ٝr�=mlYc�C5 ϛ���;Ozr%��˨O��}=	@Y��S����xz�-����j7|6d�Β4�'���[�g�-�����x<��-`�z��l���$�yXR��%�PSyQ�'Qp��Q_!x�'mˏܥ�]�7�3��uf�;i�̴du�D�#��cYQ-��F����<߅��UD����j����)%3[��P�r����ip��,�w&$�N�I��W�G*k��p�0Ǭ1�vԉё�	Q�/`��>����ѹW 6�K�_k���`*,�'��OȦ��t�/7��$���`�؍R13N�L�,��|�g���<����l��s��3sS~T~GA-
��>,W#�������'�U���-z��ǂ���sе(�7,/:����l���b�2?��b/����W��R�������Gw	��E�S8U.���@+�  n�
��̼�^h�7�P�qvʺ�ڞ�#�7:�9_�k�_�@����r�XƩ�Y��G�|�-�X~-��ӝ�Z�՚戴�N�<���Ƶ�'Y-÷�X�U,��M�kx�-��:�i�w��B�n���q�c� ����Fd.-4�h�S�MT1�C�p+<�*��lo.�'��"'�-�� Aъ���
Ōis;��]��#�d~I6o��ƺV�c��[���`��E�-B|�e��/�F�f�>�|/e]�t�"$����Y�d�:�g/��h� ��a8��4�bO���WQ����6��B�Ɋ��C]�A%��%EV+�Jţ|$�8�s/��h�(*�{����[+y�Hu��/,�r
Ap�L�+Fh���(�;�+�o�նfXd-�م{�0���-~xJ�����a������Inʇ�����mܫ*�)�2ٔ�;B�9�ܝ��I��s�G[;�.��2�����)�b��c�Q�^��U�0*_�r�m��U�nCz< ���/��퐶7��� �<􊲔�V,��ʏ��D����D���Z�)�
���Ǽ�)���M `t�Z�+���I�����]vx���#�lD��������Vý��>֓.�3���kKl8�>� ��d��uԢ���7���g�R��#x���Ru$��g�����drQ�b\�m�v�LR�C�%�| U�)��������s�SeV�i���z����+z���[6��_�4`�~�ɒ�"��쓱Eo.7����O�*��F�����c���S@X�� �c����r�E���C� ^�/Р�cq �b��� xef%�ba%���
�u8��U�{����2n?��x���Y��*����#��s��[z`���ͽs�D�����>{,�Qײ}"�^�����ye��)Ķ�;�\Q���b4��?쩍A����k��,�dz�?�Oe�]}ɤ|3��R���VT�7��`>��E(Xk��=Xb����Rz#�29)�������֊��#��V[Z7p��,�A�9B_K���c"��t�!*o�6�.���y`u����ͩ!��}_�6Y��O��s���V��\����)_ˋy�������.Z��q�R&0Dy柢a�x@PwT}���*�V6�$�dr��eB����a��:�Q����.��[�:(��ߔ�����|K�u'io�J�-kى�e��>�y��4���Ӌr���"C�݂�_M��Q�@�T�8�J�2R�x��tF��AP2	������/#6�H�uL�%N��M���|�U��E��;5Ӥ%|k�X��?��O�T��!�R�f�7H �}��U�I'�_vG(l�Y~�A_�A�T�׌Im��c�m�}�A_˿�:�D���O����^eD�GDƷ��)����<n��'�?�q�xR�%������&$a�1_ۆs�� �$�^��KZ>���t�҂��\�ӵ�kU��H��T-�:(H}��$w���h3�|��5���<�g�-y��	Gy�ZW�ķdR�L�H|��Dut�iq:��k�B���w�I��5@Wn�$5�����BU�;���>�B/9b�?̖�n��*q�Y��NnQi;�I��6S�����2�����`{�W*0��m�|0�r�z��g�l�f�(Bbj�T�A����+�v[��ˌ<ݭK]l���-�]�O����>�,��¦`i^�(����������N�Vܯ=?˓�K�-Ko�=KLr�L*qr�r�Hwٓ��I|�����r���ZZr
O�3�X=��	s��o�ӈ�\J�-I3R�?�e��]���ׇ�E�L|���K�X��p�7�;�:�?�����7�oQ�[�b��"̡�ҡ�>���U���Y��� !t�SeSjbJP>�Y~��%����,|m�чxe��Rd�Y�Ƴ}��q8T�@A�z�)�`�/��DU��� xX܇R� c�Q,Y�0Ɣ���s���*�a�j��~l��,������B��e\9o�`����8#�����5ZQV@��Y��Wgf<��X
b��,�L�\��^]o��[���]zM5Y`����F�L��D��埶�)�6���7a������]��=����1�~���@#�e*=86.�Q
��Bm=�:��YwtP�hGWJ��A�>#�p(J=�W[�w#{��X���%T z��E��'م��ά��>%?-
{S#�;�3�}��@�5�yؖ���4�)5�Y�}5�?찄@O�e��4�̅�1�plRrH'�!���A�P��\P6��<eNr��������y��xi:��T�v�ؿ�Q �ذ!�.,U���ھG��I�ј�|���6{�()�-H,AF�?v��@AzxS�oN���BV����_�/���z~�J8�QWz��"�C˯ĚĴ`��4l֣u�["�9dv6�Ru_j����-��H��q��?`�	�9�`�����[B�ݧz͐H޿�Щ��W�7�����h^f��J�1 ���W�k �j�7ϸ�:�Ј��2SG��\��f�.쳟�8l��1����>�[�s�!��|�����tV$E�����%�e��(���)h���>�1���0u��O9?+Tx�Rm檇p�hg�9f��-�*S{P�7�;���ό�^�b�L��[�z�0��	�VVڰ��H�Vb�w8�����{��?��H�;\�]�� q07��l5�dQ�&����P.倍iB�F��}^�L�:L6��7����2iw?uzܺ�z!��T}a]�
�!굝bۋ�$�F,H�u�$����BXz{	�ߥN-+ؿj �dH�
���W���%�~�bY����>ah}�:�L3顈,p{���!�R�A�ã����"� ��t�y!����`��n��Mǆ'�����1��C�V�I��P�D���,ܢ0���[%�G�U���ܘ{n�Jd����I㺪UDP�[�\h���,q_W���hy�	��I��a:T���K��h��h�i[�/�x�o�%��} !�?�j�d!���T���Ru�{���:���h�
��o�#�/C���C�!�{�c;���}l�cC�%\�M@�by��b�!FZ+���&��
l������l(©y�P0��[�E$��Qk}E��[����K���a�V
�Ώ�$hG2�e�{#��6�k}N��2�q?/��*�����X�������b\N��R�]���y�Oo�GoǕ�>��E�vDH?b6�D4�K4?ߡ�8����1s~�X�ډ��`�/��p��]��I;����H�%��(~�48��r��-����}~D�@�&��T,}h~/�&�,�}3?F���SÎ],$��@�E�
�v*�&��WѤ�V�=����-X��1�~�>�&J�av^DL�l:F"�/��t^k��սm��k�7�8 �.�]�Kh�C4E�c���+�b�?o���s{�����Dť�g����UJ�غ���fp�h	��Q^�n*ŉ���ט���z��c� �VJ����x�g/����j}�Tz������a>���@�(..c�
-�Q?eO���D�5p�
�E�{Ԕl�|��ז�+1�����`���g(,�a7�ڮ/��e�|G�,l�=�0t���C��s�$:(�~Y���-t��s���7�C�+��0t��!\6s}:G���|Zү÷�b*T~{��{e�µ���3T=KP-�>EGRq�����r���mZ��p6${�{�QkJ�7ϝ�^i���Z�O�XH�^��8+�_��G���Eï��Y������JcLW�ߎ�O"���&��c�bJ-�4�����:g$?�7�M4��2UDds���(�SX�ctC��1b�}`æ���U�(ͪĕ�6��� $��j^���@�����2�������|�'�T�l�M;�Qt����5H�!������;��f'�S4�!��&��ɓ��%#h�r։3De�8l��H���R�]Ӫ����.�|�5:\SL`�1�~�쨠�U.�TH�MZ�b���{��Y���E��I�%����«2��Ǜ������@��,���T�c��2C��@둝>�t~��Tg�]J,8r^%+8��Y������cƹ�� ꥭ1����)jg��ޑD�P߰�sÅ�D<JhSg�a%M;G��I k�]C&�z���h?�.Ի����\�5���z��xB�-b~�5�<�_�Ym�ř�����I��`�j��8G�*�7������J��M�Ju']��4�r��"��	@�b��h�?�����[N���Іr4�G��"[�;w�ᑫY�}R� �H�`[�ɺ	t>w��0����!�A�h�JW�4�/�o�Z���O�皔D'"񮓣�F�4�J|���&I]c��k�����q������0�/.v�>��N��}֡;�1�w4d���|��Y��"}S�aSv��J��&X&�#�L�r����K$�kƢ�#\�] ��S<=��>s^��]=�MQe���
�,1A��9��S�M��C[�?d�"�.�
�2\��R%K��uq��������ư�@F�s�Md�*����Vg����3�7��rw��1a��A��F��\��T�h�k����cd҇����Ϊ� �s<`?.O�����7C-�#��9�'3�L��N�"�P"�-Z�*�U��x:E�$B��S��1�U�*W `�s�lP����[?&�2_Ŷ��Eq~a�U��	s�Wb��� ���9�L�'�u�`} �2���չq��Mm
���r{����8�ȉVm���ε*�6�m%����{�2�!iBB�B�˕�����<_����@K_�O!�ٺ ��1oDV��)�� ��a��<o�2&p[ӷ����L���U����ы���@��I��
����qI���n������I�U�����s��l!�2�7ϥҽ��m,�îCI?�,ْ��IQq
m���P0�����S��8k�~��#7�pOr�R�\.���[��%��#��{���|(�"@��Zt��+.bW�9�Ij1��.=q��°qi��H�X�i��B��}6�yu���%���Z�A�.B*���QR�GhŁ��R=څ�8l<����v�ZzQ|�/RDIU������
Mv"w��C��N��@ ��O���Z���c�wI����HC�݂�' ��	�=F��<��ޢ2ʓPʈ�����ճZ���w�����M6���SP,�R
e3�U}a���m$J�H;�W�L`@���g�e6���� "#a��=�),�@:�4�J�d���=�r���1yG�K!�&�Z�;yn��d��	@ݧƗ_^J��[���f�s����
8��3fo����B�R��,\���JY�d��8F
�E�pT;f� ��tiR�K���E�d?��3�>%�m�`j0��>���đ���1z]��g늩�`>��;�I
�Ȍb�G����۟VUH��O�}�;6Z̴+c˶U�)�@9�A�ꖦ�l��
�t�D��M��)��������㱙�P�Rqvղ�����?i�o}�]ߝ��a$�.�u��E̿W��X~��ߑ
{O��'*ѝ����2�o��˷uíoڠ���ת�P�Y����zH����"�����'<�������u�8�^p�㘃�O[�Ĕ<��<���c�YJ�#HA���>��(�1�>Ni�ăD�"
��#�Wq.AFb�w��w�m�pVަK0ˣ,?(�KF�W%�Ovل�ڼH&s���z.�ֱ�<~� ��0��d��=J�ɐ$����߂�7�{g��*N�p�(���cr���v'�cJ!q��{�p���K�j�N��>X��*^X��y��	ϋ����SeK�$��:�"�*�f|=��,��a�z/�3^i$����흩a2�՛��l�i�c����K��< ��F}Hl��6z}��~��ѝ���*��>%��x��dh��a� ���������F�L4��
��V�c8`NaC����kn4ڨ����v�kR/Ԉ��U��L�7�ݢF��d䟀�x
��줯���1��<	!��������������+����=? hu���)��O�}n#%����5��6�VE�^���@��yb�]��A.deX*����|�������z���l�.�9��	�04{k�X��醬�n�MҪ��IlY�|![�����HA@�B��줳����͘Չ���m�����u��Zz4%נ?�S��C���~�}>E��|��?9x���tՄ�	G'��}�<�a�d��*�u��;�������|c�+��sHx�����N�2�
����+�ф�8�&S���N�-�#��:w(8:Z�����m��\��|W Ɖ�)|V~�pf�]W�vr\)��0X�g@l�
ݦZ>�I7+Ϳg�2ܩ�23UQ����z�퇕�'<����CU�y6���ăx�+��ߦ�0��X����t�/�F9�Vi�*|��#��D֤� �,Je��U^��t���\�.�c3�u�'�`��Ux���6�9 �A��9dv)��p@��O�&����͟���!-��˔�1���B��]����yd�}D2&le�φG^\�_�Uʀ�Z���5��=���}�F���4����3p�Q�3`��/�t�릳��%q$6���0���W�=�@6i�6���g����*�����[>�ӽ|�;HZټz2*�|j���njn�)Y�J9�`}�S��~��Y|��qժ��7t��n �c�>�OsYH;l/f31��>�.«����X5�T�e�@�w���0cT��̌Qg��l<U�b�$�8�@��l�����3���R�9 �Z(50�g�'I9����S1��F@�g�>|��b��@p���]&.ZT�CĜ
��o��r�>W��̾^5
;�<"�󸈔�aa:���L�9����b�2���N�$���;����9\\Am���4�(�sA����x���� g.���h}z��X�Їۆ@�)�:C�c�ۓ���!n��4;Ǥ-�%�B��=,�#Ɉ�4h��������c��M0��xbEH2�a��_4�sX۴�s���g��:��:�EuRKs�630����� �# �Z������?�,�2R�a�j�ձK��g��=^�)&���B���W�+.S���R[l�	mR�(z�k��B�r��wh�ujǙ����b*���aD
�KZtc��֮?s���2��;vV�=,(�Dk�9��8��� �[���b0E��$��Z
�u	/w�KZ�k���_��fj}�>�J�D������7��I��u�tᕪP���O7h�Q��hý��ն[�M��p�O  u��4����su�\61��n�q�!' ��Zqa�2-J�W&"�Vo������.O?l���11�s=���f��[�`��J�9����.��^]��d�\"G�/����N2-�ר<�X ��}
�C����-�s����k;#� >��3p��3b��cs,��1���R�& bn;�*�JQ2��Ӵ�W�D9�R$p��uq�I �Gj��m��q�f�e���f�Zar���c�|ێ��lp�r5�*g��0IKŵlm���ڍ�&ks@�.C�rG[���j�[,pH�B����ԝ��k^���4 �蹏�k���uJ���7Y�/:.��+�0��3�bL$���
�y�����~��T���MgO>n�2�g���9D�WpP�Qd��9Nnq�����e�N�֦�]CI.V��{0,�걔�'L��ݮ?�̄C^���K?����Aɏ�G���('KvI��92� 6f�Qhۋ[1�|�������w��# >�ى�Z�Ҏw}��r���hs���M�9�o��e(��|�$V����(���Ʒ	5qV�~����6sG�cAß�M�\��j\}�iΛ=)Y1��L���ɘ�M�8�)���iޯY�xPb�TKY:U���%���7S=����Lg��'���HЛAF>�n���U]�dY�r�M����|-#�H�\�H�2�A(��j
vQR,�zO0QC���d��Lp ��(C� [g�Y��]H��E'K�̒��e�TA�5&';�IQ�
r���������笡�%�^��#Ec��Ɗ����q�R�<U���= �:�q��Ft2��f�ĝ9k�a��'����ȅ��DPXD�tU<�naf���{���P̽?+�D�	:��f�|q�����+1E��1�	��BQd�#`��Lv��˒vʋܶ��¿I��<�^��kO)��h�9$���|HH}�	ބB.ڹ�2�-Ծ��p|K�e�_S��L$���8:�����ë�h�V�vT��Q���k�W�Ƃ�ȊK��o;���X�{��_�������h�ڛ�\�ş\ڑ�	�c�j�ך�Zg���O�h:j�GӚ5�]��;a�H`d���o�T�670�	4v��U�6��:}��OL�{UB |�[�5�]�����]G��,�b��xP�!�g�Y�WnK렟�,���u��N�y0c��������j
Ԗ���ݘQ�Up�0�cYM�}�fP�s]r�����*�)�9�,!, )s]��dDRo�@{�GԞb��g��Vi�ysR*����AJ�;<�8��>�4� ��b��M�e2�5@���)��k��I`��I���%�KM��<�l��mhe�������a�����7 lq��(�7:B�u��=+Fd���U�59l�8��� ZZ0�J���X�*|v��n�dI�Έa6���Iũ{�=�l�{|����0����20�2�8v��Ք;H�ے����Ŭ:���R+��'42�n�-�0O�j��Ǳ��;�����ϣ�P^q^�1~=Jڸ�?�}���<�}�'lރ��0�l7[nwj�rs	����,�>��QAAG��l2��a� �>�(J� �F{���(}�5�/ۑ��f&�)}٨=������5�)ܶ\V�7)ȝ�=�s�{CU?�J96�ZD;+ށ��V�r�:țv��zlZ�N"��@O������q�xb�5��T1��*tG��Ȗ=Cs�����m4�R�#�\��e4^]�5��{�x��Iڈ{������y�TJ�����*İ"�}���},OqC�u��X�"%�o�I���G_�6�H)�QvȞhʚ�_n�=M���jwNǦR���Y؞�������ɾ\���-Ʌ܍�4�L��wne�r*s�2�%�����ɬ�%�Y����k|���dOv���B���nQ��{��\t5\�������~��j�3���ݎ�I�c6�?L��o��Щ���v�N �%�\^/��qE�1c��_N1�#|fY	�6tbއp��VSߧ݈���Ӛ�LB�KJ�!ͯ��>��{u�(����f�ۣ3P�T�t4,t%�"I��t��M����Q��]3���~|��/\Qw�:�ѵ^e}���?!�
;�
l�|�����Gy�-^��ǡ�P�m�A��!��(�P�I� �6��:�Cl.Bh�n�45UWx���ߍ�4Vk��#���hI�����
�7��g�#��j L��P�����L������$��V�P�&��O*\vۓ�D��L�qUgMq�mV��@vQ�s�r?�.�s'�]5głZA�7�䪊oZ;ݕ�TLmh���(������5�g��vݱ��ɣ�d�2T$�b�8^��jI�����V�[%)'����u�׸|f�#|��0��c9[�Y[�(��<U�a�C�I4��n��ի$Û���IK��􂗮I�ۚ��*]�p��"�4v� �F�ݶ[]<4~�h%a!�H�b��=)����)�aY�wv\���#ۊ�;�#S�~�,ǌ�[`�]�26��2�Ym�8JM����: H����	�!	����%���LPK8 !���u�a�'����x^O�:�%��\[`y�w����Z�K���e����J��
��xm��MC�Z��oQ��C��?1G�{�GD�ʝS��ߵ��U2l���M���c�Z5�2j�:�*�ţ$��@��EC~�n��R�ι�=����X�F}`� b>fzU�]�Hv�[�ݢy�'��W�7|��P
L�-��@l@0Q%�s��f-�h%alx�!I�T���m���Jܬ��g��&t-m�EY�@0����9��ϸ�3CC���=�Q�z�4�e^Ь��~�����H�ȟ\+�����|�D�����*)+�^^n�L���Ӵ��[@'����l���|,�܅͐���;���>�k���5�)�:�t
}��'�����g���E��~����`s!ĵ����X��J��0_Yt���aM�5��9s�P�df�fb�����~D�V�����o$��$�q�$$��E�s�,Lh��O�&�SϪ����{u.W�8dD�&v��ڸ�5�
D�5�hBf���	��9\��Q�Ѧ�1.y��D��Wߐ_��Yѕ��Tg�O�Q÷"ڐ�������ɷ4������6҆���Y�g>�G�RӤ�JO�j؆^>�������K@����9
z�̜f�b�Ηzs=�r�� ��IalW���F��~��b�'���`:J��G�G�!t�c+�Xmti:����Pr���G2�"��%K�P��e�G�n���%�K}����n�ʫa'�y�u}#���������D�Ta�	 ��셎��l��ܜW�C*�?�ܟ���yQY�C�Y�ā}���;���ܮR�*o�3�$G��W��0r�pT�
:w)��{��i�Gat�a79��x"�@�_\�O1W[�l/�X�h�|ٌ�p�c[,"ۉ�6��v{�6�&I��I[��X�j������.ѿ$WD@�v=�H�!*]��+H��G��� ��`�F	�2��3����v��u�������"�F=�pC�6g��P��L���r������ܜ�ivF�--1nxt;h,�s
��2�*�B�[	���"ҙ�FN�Q��6�p�b����AS$�jP'�)X�D�֦jjg��`oTw�2�	3sbCZ}�e�M��%F?NO�J(�i�3�j��cV�`�Ei)\bw�|u^¸��AV���F)�R�>��p�E��0�'��¦�@�m��l1��hܔ8(w����_��\;Y��x���m��C���&ؾa�z������ȱ��i�'�����&js����)(�,G����hg���B��i�WQ��2�e��+���/͉տ�fQ$�E����-�릵� �NԶ�uy5qT��RrR���A�^�e3dbU�)�BF�Ɂ�����x��e=W�[O6�� �LU�QmR��r�$h�&�9�?��#�ց�9��.
-ًB�%艕���ɇ�mȈZ858m-�<^�c!�[��y��+�;3�ْ8�b�ht�\��w�&����۲_ȔX�A��5� 
��$'l"3[��r�)��2R�ޛ�Nj+MQZ9Nґ���BQ�f�K�p���'�ӝ��].5����Qâ��B���j�n���H6N�]���M�P��b���=I'��a���e�Sj�ĀGX~���Ӌ�s�@�,�*C�K��z�Ö�mgQ⑹�0ա�S�h#ڐG':����a哚*I�׎�	֪<�5Z]�D��-.�=?��b�� j/` M䏽���H�7�vS:�f�-�Z,=���v���A͸�P\�`FTPTNn$зw"�/�����i���@��l�0� B9�[\Py�]4:�i��\�7�h�.o脶�P�L���t��ڤ��s����c`��p��I���l�K�PK�\�գ�='��W�r朡��u��!n�B{�Y�̆��u����]�a|bR�҅y~0YZ��hh����3�	�%5�pӧ�\[[69W��� j�wҐ?&x_��5��cc�s/ݹ%U�ߓh9y�<ʶ�N^C{�蓦��XP��:Ϊ�_�&>A���z�����,Hu���������n�A��@���@U�9vw?n�+�9(|�Ѣ]"wD�h%I��D�9��^�Za�6�%�ڊ�[���@Ewc��~~C��m4M�H��N�	CQ\�N�o�e9q�Κ�E!e3
����%A�ܸ
H��u�E�@J�'�}jIˌ�v'�f7� �����P�UbU1�^���H�Z��Oe�M��x6jG�Kl���bQ
�*h�u=az=� ݺ�wI��i���:0ݹC �7�	�(��N&�����-�H�-��������*�r��i������;��ņ&�4]Ȑ�L^;π��B+q?��HN,�j���'����A�#@�No�>�}K�0����N*�wED'�Hc� U�P��εl̈�ڼ�Ve{��<�@a��8��O�Ņ�!�yY�N�އ<��Zy>Gŀ���`w�4:��x~�¨��YP���' ��m�Մ����*e� �����IH��{Ϝ)�����<����~&�D��8�wK�^�/8��a��D��zU8�^��ș��{$#���s-1:�����gJrr7c�Z��oO�qw��-���H��Դ���C����*���I�� &��P#�A���D�$1ī�Ĳ���_�7矺D'P  �������=^!Nb�z�]��bݞS�L�*�N�\�F3�`���[�b�]��p_=�*$H��� vm��c�k�`�<�E 6G�L@P�"�|�J���t�[�񖨜��f��` `�$ә�.>P'vfkg�U|\W����tWUֻKX��$�Gʧv���e�Vq��X���+�Lo�o��i��OfD��t
�fb��O�v��q�1:Q���]ak?�q�8Tˑ��V�rU���}�y+�����\�N�;�8w�������\�M����qc����J_;[۠��A-_w�ф�w�Ћ�-�a����x�3x0bT��7���[	��vI�}���Jg̅U�dL
�Fq\b�i8�����T���i^�65(������Lf��ba!a9zX^̨3�iAڂc�VG#8X�&y �����i.��N~���D���T$�x��<G �w؋�r�
C�n�]�Hy��=����?F�o0�����r�<:��6��fw6v��Ք�o�io����H*`<�8�n]m|n��K7���? t���H���3�(/S���Z
�u[��)�U�� Џ)��c��pҧ��bB}`�!DG
aJ/dB�-��o�P%��������N�/�J�«��Z{Oa8]��:����y\N���E*���.���l�?R�U�
XOn�`s���x
F������PH&%�l$N 9D�ag'��N�ל�)�E���_�����w#���e�A(�p�n��w���F-$�j���vVI]����n�j#%!�0�=^��4VɅ'�"�"qoW⮀�?�V���������`� J��U�5)�Cpj��g	����rZ���n����
X|�{O2��U[@V����g�����$~Y/�f������6k])���*`v���L�Z�2��� G�2��C����Iձ?w�Pk��T��W��y���0�cI���<H2+W�J��}I�4�޸2� ���Ԍ�<Z�d������(ԧ���%�] TJ���%x=Dt��T����cIM�+9�τZg�<�;I��?m$����	�g[�xv�[���
���ծ�:�i$HV�࿹;�F!i�r���z�$�qG5vq���R�NY�u�}���a�y��pe���.H������||!�������yxDkx�k[��?25�+ö�WΥb�S<�&[Co$���]-�g@y\r\e C����2�S���e�hJE�t���1s�"�uo�e��Ïu�,�Վ>}.	ry���GN�	Ib�#9A4h���[���>F�p��J�a�#�xD����q�x�^�Ӯ��tx��@�@P������ݳ��|4�=�ۨV��N�i�p����$�=U���j�Z����u�� �p��%*[<m�إ��J��L�4SOk�Zt4��6�MDY�����c<?��2��pa\�??'S;�G��H�L%U=���1�<�r����oq�j�
�9��5ɫ��Ll%յ�d��zRt�ر/�R���x�D0�h�M(nf�{�r��z�K��\:���ZwQ�P@�d̿�bpJ
J�}��s��M�jk�L���%�6�>��0EF�\��븆K:�X#�9�n�
ID��q2`ʖj�(� ��$j:�=�z�n��vY'�Q-b.��ْ�t�l2��W�tmEJ�ΰ�!��hax���8y�/S(ڂE��o��s�@V���||�m���G!S]h+sP�	N;ߠ�^X�	)����}ܥ�A�F�c��t-5 ����Y�B(lX����@������螧|+ƭ��B�{
74X��%G{�)*��P}}�a;���������3Ă�/�(�l�`�g��|@!��퍧���
`���S�|ϦU_�f�X)�)��į@�x*�K��U��`P��~��`0c�s�;��=����u�6�G������F�t�"ݭ뫋,:	$e`�Ș��CuI2����cj!f�/�hL�t-D���8�J�UN�� ��+:�$�&1E9 ��,v�Ƨ��1�̣�d",Vz%�	�BV,=w��qư�����z���;ް	KK�b����M!�s~�H�9m�,����Gq�ݬ�䏷�ta���.w�i���;����;�"�(�S跟&*�+T'����'���
�K�o����Ե���{9^�(:z�,ᙃ�<Y�y8�'�L������ ��N�i7�fJϐ���5u��1<�/����M�|�f-�����wQQ�+�g~3	.�V7��n�)}Q޶��>���\����!C4
�	0.�Ew[����^�yޒ\����p��R�R�Z�@��{ˮ��u��3�n<Рx����.��p�ȅ��.�ۘx~�g�A��6t�-a4L��n�Kb; ~)J1����Y��ҡO�)�iuҢ��ϩd#m6J���n���Es�t��	֫�T�0�����a��Q�Q���4n��4\C+�F�� B�l���S��]AU�)|�3B="_�T�E��o�zW�4r�k~�X= \����ז�KG{'��i�~�O��6�ӘX�k���+p}�1������b)/��όYt�!�0Mzz	{C����;5�8���؈��N�v�gzD�����fVY����K�
ū���(��\�(F>G^�/�A�/��K
f�B,���&��ɜ�2�7S(y���}��}�X����K�����I0Y�8`y���C�HI��o��2h�����bpaX��|$Rء
��C�lR0��
�h��bj ��}@�l��d$����7����X6��0�h�x�" 3��=p�0 j�������&�ɽel��s~.0��ܒ	k���{��K{yV�1��l>���4�~�N�[�ϝ\@���Z���L?2�O�9_���n�7v�� �u����̓4}�H+W�c�6,��ҫ��qi�@�9�wh�J�n:���!y�F5���	���������������Y�7.��Q��L�N�h5��J�2�L}X	�b�)�S�M6�#)�6�m���v�.Vx��~�I�$�=PT2�1��.+ʂ���;�mǒ����v7�a:Q�l�j���B<�FinF\�_���S���u�ᖊ���]�팁���o%�����9<�{b{.BU�����g�!M�nh�������hK��ɯ<3�,c����X�ٻ�~�eE�#�N���S���ٱidc�M��!���w�6į���Ņc�ܗ��� O_r(}�pv/a��YQ�}�4�L4����f!1�Pc��S��K��!"���|,]&o�חa;���*�^hm1�pt�)`�z��o��i �0�������Wv8ܱߕ̼H0C����3��<�)n%��L
V�B�#����sf^� .����V�������Ӕc1�?mԚ**q��}X��Sk7*�#�-�N��>���$!��8>���h'~��ɔ*�}f�F�0��j��� 5#H�AJ�"TF���K�9}������m^o͉e}8d�!��A��Uuu�Y0i>1�޹���1�S$ɖ���>��f���{Lx�Cr�1|`��Ԃ�7�j+�d=Q�Ql=�<�3Y���]fYG+�k3l���+����	��e��-?ʁ�l��b���8/����G�8P��j=t~rJ����>�]f^�"�� l�Vfxk�#�唙s�9w"��=Y���F
�g��^�i�z�>�D� ���oj�ָB���j 8�̌ueᢋ��#�E�Yx�Wr,�Nr����7H3�C���{�H�'T�&"w��%��[5;�,��KvE�^�M��̋�~��*9Ih�L��)O����o�b-}K�hS��oIL� �!yւӿ��[���w5�KOl��&�aLA7�uE"��f(�By�I�ȴ��5R򁨓��B�BMM���k�8EX>���!���!��O���;>����Ps�s���6����A�zϽ>86΋H\y�W�֤�>tg�f1�,�6�����Rt�nԊ+������!X��;`)c.O������D�ȡs׿]�X��[�"��,Z6�7�r�eB�J{�����GPM����{���+t`�0�{�[�.Z	8�-��)��V<	��m4P�	��%�,/��V*���:Oo�=���_���Į�Y�����!kk�������A��|}vDo�N��B��|9c�B�M8	ש�,���>���<��P�h(����NӀ�����v�A�k�;Ͱ�sq�k�f t��'yN�����{���dE�*	W��G���z��k���,�e��@X@���g�^�,ŲTΫĸ�Ej��6���4WD�}��@Lw���6���A��� ]�J�bUխ���Ǐb�3?� ����9*O���b���Лt�9����w컑���HԤ� ׻��Bq�i���[3��eDބ[�3 �
��G�_Q��㶍T��2���5��*0�A�b�I�g7�GP�WDBtՇsS���"��g�D�(Ov�?�#uXLm�`,��XT��1���� ��i�w�uw�Z[WPK�KÙT�gVw�Q����s�l�o���!2~��Q�����X�~U��q�� ��`��vv��	㤕�����(��Y�(1�]l���_,%������{��r���:iL䔼^.����H���<`��j�ֶz�d�>O�(�"���8��R.�Ii��⳽��)���&۴�$x!;N IX�}Vyp臺��+�)�����|c� ���L�鿮ߊ��:;��ߓ�T{q	���ZZEw�� c��Ȗ�0��	�#q\�X�#h{hI�Ƶ�<�`LdK�������z�]�[:@ϯ��O�P�J/l{=P_��\�UO���7�-K,<���.C�Fu���f+�P�F}�����ွ�Dpd�y�
dZ;�^C�|0i���T��C�~=�*P���Y��M#z�m�㤭OIn�o)ɭdV9xRr�h�Ö��^viʍ�-4I�C��Rl!W�ڔ�1�a���58�7\��ј7"Q�;~�z���?3����Ģ�ʜ�����D����YޚXt�Oґ/Ú=bDʑM���>M�g�C���������З7f1Mul�06`��;��K9I�SswA���Ki31	���k�g�p�۟S�'�Y+: ��@ګ[QM�_��9͔���O��mS��i�����F��������;Axj�v:�b�\eP�Q�LK9�,♜&bm��Uj����j���͹�νKv*��8�x�PQy���]ej�n���1��D2g��S
�]��0�檻���^�Da��c��O�j_#}���	=tm<{?�¦/�]�L��;Ί�}$Z���x0Z�N�G�TA{�=�I[���� �l�ٕ*���L��64�$����`�lI)1��<��zG`K��$ȕ|��ؗR�Ŷ��aǊ�O�o�����-��E�j��!�� �l*����8Ym�G��v�o��P���{f𰷦�c1�i������&B��m�54�����M�>8���l>�i�ݽ�H��d�U��x�{��8�� !-��c��d�䷘����!�U��Ʌt��h���"Ս}!�w�G`�݃C�[�Oi?�����KRF*T�-R�	�K�V�iH���,>e�yZOӜoҫ�.�N��)�.�  ��J����c���.wAK4�G�;㾋$��3ޤ��-(��U7��(^!@.ʐ0g��w6.���(�UWΘJ����Nq/5 x4eY��(��&2WO\�f��}@����$��5=Xv��(���b�DF3�<'�80���T�MD6�����o4���[�1v+od]
��(������>�T0|����&Gki���ҙ���P[)�У\cC��C�4��D�M%�[���ga	]&͎n�MF0��}	�[q�Mar`6�����C܏�|Py6O��$IV�ކj��Zd'~-4��/O��B������L�������lX
3��M�0}��AX/�\���n���=�Nހ�-�Z�EAr��UR��*w��PA}��ӵ��9�o-a�0
��m�]L��x��E�S��|D:��B�O���6Q�n�X��پKdY�z�G�p_E��Mru]Ow�a?jX�K�X�b�7ikZ��	Zw� ]��F"�K5R�+ȃW$A�W�:Yז�3Pf�:}v�Gz^I*�CZ/�K�v��
�P�Ɉ�U	C
琠	��5'EG���ˏV����b9��E�yh��^�{����,�e�����M�O`�}��49�|S����A a/+*�|�;����B��i����p��7w�ʱ��-8'r������Y�[c��X$5��=�ó��;��'�&z��K�CT7��x���hx9�,^�����+���?�0ܱ`��ҟ�,$Z�H:�=Z��c����c�:4�/���ϸǳk'7�������R�s�|����v2B�V��p�L�n<�Of���Di�/eELY#��,Ts�����4y�1���=�C������kw���#�Tr�Ex�-�̙;� E&��c���cm�K�5�-���jH�7�1��r�{�hð/�n�L�/��4���m/��Q�mu�La�=�'�q��@+Q�:xb�ϣ��t/!Q�køDz�/�㍓�V�n���>AB�����z�,?E���*��,LI�/��ilZZ6�����X:������P�k�.�B92oh� �g h0�|���|��:�Ę�\�����y�ʝ�������
��{UN��Zz1���w����MP>$Xv���L&����q�Z��_	,yf~Z��޺�ZR�Z�>�@v�Gf�#�}��͑����Y�H
�̍`e�h8<B7Ug��RW����B���>�G�4������kf���G9�e�{T��8��:-_4^��
��ݵ�q�S2ɦ,!c�4ޯ{��wQ]��Rk����8SM=v7[��O�as�"���RCt�at�7�ߘ�1�]�	:恼�O����&"WƧWh���9��`��嗑�_U�6e�������3��H<�MBTͅ�c�pl4�RX�����R��w�C�f><d��d�v3k�%�N@� �2w@�wo��;s&���*�&�F�C׫��9��_#E���_%V�������)+ҵ�x�\��۔����x١ �ǽ,p�\�*e��Ae験���ձvΐ�yrb{��K�#���G�o���Q��r�f������ �U�_�o6����i�L��ď���[kM�{�k!�6�f�B�N?�ʁ�ǣ��-��L��N�V�uK]u�w}�����Rcrf��C|���Vܫ�7'T�i�+���]E � o�7�~t��a���$��eF��J,���C�xB��l�q|<=*n����c��t �'�UrQ�7�ShP�w���D])&7�%�Q�L�Y�4�㼔 [��*�u$X������@
6i�X���)�F|�^�!�u���|XD����چ=zB�`�0�G�?��1�A����0���g����
��