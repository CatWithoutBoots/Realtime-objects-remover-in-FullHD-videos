��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&r�F���oh�hi'n�į.2�-`(���ggB�]4��}�T��mJ'*m )N�_�6ն�4�C�������s��q�����Z�x��_a��?^��R�b��m��G렣���}U���N
��կ��`ڍ �BW����C�&e՛��Zu�E���[�/:_��!An�E��Hs����7��5D�.�<�.z���;�m9���S7�V
'�=Z}H)DV#F���WZh8 5C�K	�B[�@�`�U��*�$��^H����Yz����͔���L�o�,b�&<*d�Pӵi�V>�b/�J罹�����5qDg��]��X���DUF��+3~��N�	+#�Q-{C��?�VLs�	q1�6�N���龭�n(�#�Nr���d�lbu� ���W��lg�%���S�wy����z�:if6k��~F9���\��WfW�AVT�J@g��v�#p�d��͕E���ƌ���X��[�RYx����lv���3��~
��>a����l֫N�*���,�B�%5p�o,��;�?
^^��rJ��q�<<��Q��j���mQ��R�a��:2h?3��P�@�IH0���(fHG�M���ܧ�	�r1o��Sݮ���kJt�5X&���l�ڴ����"+Hu<�:�� �s��^/���<���X�#���5���v�>�b�qL[Aa*�����
��sܼ�Xwո����0#W`�$�o�2G��l[q`x������r�A��'�W&���136�����VS��%�A{3��2�4�o�]D(wW��ؓ\��[�b�w��t
�opC=���i3��8��	q�����8���L!0({����[�J��1胍W�������q��&�ǵ/n��ң�.�j���۩��Fg���gq��U�d��D�}pqk\&��vI-�2�ѓ��jrSC/��?��p�΢K+�}��b������0(L���n���NdDW�;��C���K��p��N�8�oϋb�D}�ꎒ��	�a�䭝#��Zg����ưϾ�E��C�\rd��̗�#�����7�0<��T֚}-�M"SzS�p�<D!:q˥�ȱ
ό�_+��q���Q^�4�B��g4]�&7�������М����UdUL���NT饪 ��:et�wc���f������i���~m6�#l�of�bu��Pn��%V��z�B���2��e�(�t�;!\�G34��iCJ���A�������� "������\�����'���f�J�O��V�q!�F9_ޘ�0���� 4��W�Ry샄b鎶�y|�֫��:46�"\��zK���(�����I��*�����~��'�f������d�P6����zQ=� �TG�b��NoO4�C��yw����}��9��6~�e|no�=��ƕ����,��9�唉Qu�\�~/}i��R�]J�V���!7V�h�7�/�n� �M&Ƅ���.KRK3#�P��dĆ��Q8��L��F�kz��Lߡ�5z���r�;���a ��B#�5���#yB�\��)��&��E�.kh@
L��8��Uv�R��ӌ���Jx��X�O��n���\#��[T�(p�� �W"b܏0sG[��)V�O���q�v����%v�08�Kg��M�eH�g]1�Jyv���	"���K�Q���;�G6�E3Mb/���6��)*V�j�%��V�]a��� ���D�ئ�2Ȓ��$��1/mňy!�ޙ 7 0���l��x5��i���6��ת�@6._�?�.s[%/+e�zwl�7�����`�8�/~��q�1�}�!,�O=_/��ߨ�VU�&����9�[��N����#X�|���dS>��g���u�s�z���	�c1���=�$���*u��䈂K�tXq��n����9�����'�5�Og�Ɉ����0=��e��e|�u�wG٩�%\z*�hi���a�&��I�.2�L +����b�p˦F�C�'J������
�
�Ff ?����[;��#Jj,��OY�Z��~D��y�~��	��DI�y��o˯l�:ĸ(����!A��J�/i�6
R�Sq쑳�-��ݺ
�x�$���)�����'�_�%�zt�9Α)����Q���h3�;5����n *x�d6�l��l�.�d�ϢQ9E+����<K�$�Gi\��Dc�5n��'�R�'pC7���ZpwQ��8p�Жꔗ�Њ*�;�і�FU����:�
�c)ț3�"��j����<ȱ���&�� ���Ù������g���\T�d)!�=G����'���F�wd�
�ېC`��0h�O˔!=�ش;s�o�@�̌I&�����x*U*�Ɗ���D����mi�#�ꭙ�-���k��ɫ~If���j�����Ī���,&jA���rIiR֎ԝGc�6�,Zca���E��s��
�_5D5�n�S`e�Ԕy�o�0�Z�up�'�[5�0A#�_z����O��7	��znAPQ�x2�bk�[S�e?&_��]1?q;�):RK���4Mm3v��,����H�Í���]�jkT�y�:�}G�j)p���.�i1g�'Ǔ@#��	�� �"R:۷�拱xzmC��Wi�c��$d\���0�	ȶ����9:Z��K�Q��a����������DY�|Z�D�φ<0��(�#ó���]e�ݣ�.��$�7H�T�t�J�T���y�'��Vj�p��.>V��s"��#n��g�9����$�����˖A2�,/tu8|��τ>�k1✐MR!����G��ˋ���l#�ܾX7"�����o�߮n�o�����?ٸHnM���)�����]! �����p��?꽃�Rr�QՊ\C/�N�' �a���E9�괵���X�*�ɴ���J>�٦i*�"p�dq�����>��L�bXy�0g�pOc�{]�(v���@��jV������8�L��"���RsK���{ҭ��5`ao��$�V��(�c����3��W������"��!Sw�x8c��+F��U��R��2���|Ӊ�ͻS��@� yy�jݳy ?������w,��/��-kfn{���6�.j4�ԇ_t�W���~�1������;6B�_"����~Ko����tV��l���%�=���ZTz��.��±�<S��L��x�3���r/��b�.�^���_(�x�'�i�tw�4�.���]ժ]f11��q�2
��W�B����ˉx!N�d˧�x5�B4��CO�3�Xlri7�W��ܻ�v�7:�$��u�r����n��a\����!�r��T�T l�j�,��䈷�YE�&/�x�����_B~�޸���w�������%��ej���}gƉ6����?A)�r 6a�r���	}M*H�@�տ��>�dz�A�zC���.�%����J��1�W�1����#�{ ��K|���t��%�B��Y@�i_�B9¹������}�1!gBnU��-5.z���nb=ek�}�ܱW��� ��H�2����S����ho��nb��TL��x5V�@�V�б��x$}��=�YE���C2�Ca��s6�#�xIR��(8�7��kI�ړ#���=լ&�?�T<��p�3�L��X:8ڳ�	�b��a!�����덢��i���/�4�s*�"�ίƄ�Ó�s_W��fF��$�x(ųil (��&��XT �&��`�G����s1�ūB�:Q�!��̗��7��8�<8x����X�A3�t8<K!U��V�}B)׬���ϛMАB�ȼ��mH��ɾl��%t �����-B�tC�/�i�
�<kj�/�m>��i7K���x*R��:K�5�"�E��0�z�ѻ�yY눣�+o������ǞJlۥ���|�B�;:*�u�P����r�����?��*+T�¢����p�oع�OYU�G4/H\"ַaO��au���c������$�!��M*��o}�����w,x�R@��w��%��"�ۨ;%��u�p�t�.�x��G҃��M#4�":8UJOBjy���t�E�ƻp�Z	��`2红z��pR5�rk򂦅ֹüE
�8U
�cłD ]�Za�u&�zS�hO-�AR�ʹMk��.!P���6��L��Q�ۻ���> �7��4.4?N!2m�7`���+5.`�UMu�0�6U����Tl�;�-�&y�û���R���2�g���@C\��S���~� G���*�Eg�߰�F�i)��67jܰF���T�:�(�cc�qS�O㎪[;��G��&+n6��.��B�a	����6vU6��� i���
Y� ΃��s��?�,R7c�2�����U	#ȴ����bd��[��h� @�4��Gs�	�k#�ޣC�����r��I���ݳ�t�!�덨�[�+�>qhqr	n�V%:^/y��D�U�]���f�j�ヽ<`F[��w��0��M\y��2����/����f�q="�Y���|����0�:�l9cY�2ֈ$#.P�~����x��P�����������u�h[���mz��U-�C369�qK�W�n+��>L��I�L�zC`
#��ڌ1�#.P������͚M���C%�c%��O1\v�x�x�`��GО���3��ACZ2�����M��Y|��ת��2-[��|�6ʺBz-!hږ[�S�Z�y$'�U����t�0�?���psӰ&UĶ�;\��&��d	�S�r��OT�]j�^ӭt�j���f�X,]��dp`#�,Pe�iK�E���*�Ζ��
�H���D�����(��Us�焱����=;��o���َ1�A50��eS��
�O�������������<����� Y�⎭י���B{���)��������`���
y�0�vp������1N-}��̱�g��)ѩYJ	�����.=�t�qQd	p�U�H���F�[�p�NDg-Dp�n�w�=�n�d�f��p	g���kK�q��$��ꣻ��TE�DP`�/>$;�,h9t�$3"�s�wk��v�.|_�Y���죋/����
�m���<�6�Ɖǃ}ث0�|��	Y6��E������i)�r���1�5�e`4 �E�&�R���gዂ���#ȡ^��8Ǻ|߮hX1`�.�]��oe����v�r�P�o��9�����@�$<d����w���	�twM���[���*���e�l8��A�����o���qu��?!�#R\7崏����~���c���垙=�@ ����(�<�OӘ��ӷ�Y#�~`eM���:8G'E�HM�Tg���j-���]�}'=&��!5O�[A�O�h}�)h���.������x����*)T9���&ʀ���m��V� ,�u���)��K�s��(GG`&F�Ƙ����H�M����������Z�?lS�u�=1o�W2R�h�!9{�c�!���1�T�N�Q0���wj���`*�^3҂\�~uDn��ܳYFx-X��^�"Έ�\���,�ʨ½Щ�G�0�/]�Q7�b��S��{>�Jf�6J_9����s&t�����xX�10��� ��)P�NR���������P����[_���A�oJ��t��u�z�� �Q��׸l���yD ����j.��#�����>��66��ȚO[���WU�B���H  �C9-q�� ��� 7]eF��(��5�掭�"#�����'K:����lA��;\I�y��t�ڝ������F
)�;KM���:���Ta��Pp�73�v4j\���ޖ*̄�Fv��O��Ҋ�b�U�L]"�!�'��_\����K*�S�2�A�l��YV���T�˙�I����*rQn1ݾ۾�;�,M�}q|lg:�n�����2fpj%D�aװ��~k��2X��cC�I�{M�R�<[v��~B�#�N�! k��8�l����rE��e�d3�����0Wų�03|� X�2%�cұ��Ȏ@��V�4j<���~�v4t�&�P������^Y�X�"|<h�6.l��V��m�a��f3��L�^��u)� �)&�j��{�`jAUK�m^� �Gc�3q�SJx#^�����7�MC�3*����I���3�vkȏ�QQ5�1�c�M%_pu"faԉ�WP�@���7�{ޜ���KO0���E_Ll�?I1���D�Dy�t��
���ۺWk��#�"��"h��S��<�jpUM?>����ȣ]����r'-d��7c>P%�8�$.��&a#܍����Ή�N�;�C��n'�F/�ŀ%-�P!ӏ������k�t�7*�E.����1�
@b��%;e��.Qb���P3��4|o��c���'[L+��D����"��=�[QEg2�'W�F�H���7�(^~$?�e��YkXj�%�@��/�#� �S�G�7@s�2�À��7�!�,��>ݎ7���v�͞��G�$�R��$K���ԪUފÿ}Sk�*����[�E�om�*Vh�:�1VyTn,f�2����ϳE%�����%�w�$ sr����$jP�ט� ٯK���ؑ��-.������qa1F�	C8�F=�Ŀ_��
�*bm�e7�X#ʩ�F�8�������L�G�5��_]#w�eS,�'1?��E��$��&|�GgG�Z�3����#�d]q���f�&��!wS��
f��f��kEl���b��&E�Fw{�R!l���G�&��<�YpT�\���x;v->=�t�w�`ߺ�̪�+�={������2�c�7o��HN#H��*��b|���3s��`О���/΅P��-��`�F�>$��c96�F�c�����DWa�<	����JW�<���6ET��
&2Ok��w�p=�AQ2�wK��G{�@�Q�B��N�_�q/��r��hdG8Ѧ�����cF��!�yt�Z�r���)���r������:�]��s����g���g�p��/��6]`sk~#+zv�sû
BZ�/%�}Aq��ՃƬ��(�����L�u+�W���.��ttW��W��.T�5���y1�\����Z�|?V}�=���	�!F�J�@�~�q�H{�]�����YQž��L�	�� s>QE�|�XDDj�8�;&e=}���DD
rՉ&��&����~E\JAx󉠰7C$YߛT���2
r��6���W�1�m��8�q�ْ��\�ȇ�=�~\-<̡���欘 A�L"�^x��j��+��M�{�8���>#����[ޚQ�ԲS�o&.� ^>�l����R �쥺�S�f1g�Y�Ղ��k��tz /|�b%� ��EI�-�?ܷ�G��D�}N��9��� ��o��i�S��NBJ�q�&�j�qDu=�,�SY�`�}����kK�V�##S�؇*H�(NGd�ۑPs�Դ�3��Mg΄چa�SA%٠��fn�w\Կi�H�p	dn���a77ز�`	���@E-e��V���kd�j`"$�/G"9�!�-ߑ3��7����/*��"�x�Zۂ��³�!P�}���&��X�������[ԫ��n/�>XĿJuσs�~�,K���s��P�����xW�Ի"eE�+���o�,nJ�+j0ЯQ��p��#�eVҥ	���}��-���B˃�*m��jm�r��V<��?>gi�K:��w�Pv��f��YW-R�1�e�W��2⛛���c��
���`S��|6��Di��}�
���e*��'���'B^��_��.��h9�3�q�&>n�p�@��&|ʻQ�
���4e��ɇ�Ewl&>�����D��H�)('�_����i�j!��$�����a%FD��i{���  ^/�X�e��[�V�l��m>(x�����͞���������%�+)�{�L�ڡ��-/3�ܴދ|R�'�d�J���/#��Y&�6VA�ѲP�F�r0� t����. \���L{E�O�:BЙ�S"zy$�)���h�����|��̋PX�ڞyq�ɠY�U��T�z����1m�Wn}�@�4�Ѩ`eN��:��v�JgnO���l��.�T�r�bs���NE�L�!��{��M������H�/(�t ��s�]�$,9�-�\Kqs*v]CKc�l��,�Ƹ�B���%��V&�x��HBQ�c�_���za�No��eh>�L0fo�?I���_Mb}�1<�H�{�ܙ��ʼf2�Nm��0�X}_����z�F�"] ʤ8�XoɇWNc�&4�G����^��H��G�j�}_憘�������E���"�F
	)y/7���3��y�"�ڣ�F�VF�d�K��,����<��b�۪�������|vg�Y�U�{����//����;Z�h6�{�75�Vb�(��B̷�y�ٲ
���<� #��P�e7<�.ȒX$$�3��B���_=�`0�Cp�%����?�Ec�J�"헏#3#>(\׹��+2B�d��P�����k�A��]'n"�ϙ���4:n�f�d'v��̝�rK��o-,��<[p��v��L>���x�f��&��O��G8}�*�n����@�U�;�O��Pn*�.�/;N��؜"ji���i��h��E��9x��.�rg�x����`�
�'$�p���	��Ji��+G�W4]C�F��j�|{�ב���4:�O�ж H����T�G%��u`W�]d�$���6f_U�Qy��!�E��(��J�'��NI�i`��)[d�����M���-<�ep����?A�=�κn���9�V*�?3X��L����(��x.?��D��OE�<]�>]��xX�#���<ԦV�©E�#��7�sC�<<��)~��p��H�� ��ex�B�����rwVq�1M�_Q��������$K�9Σ|�rӬ�=����&�+��YmW=����[D路2Q�R�t�F�0o���B�C�^3E� Q q��T��Ot򅯳�$�X�'^��-��kRr�jW��.]�Ng��C�A�	;���R��NXW����ua�,�ߴ���fs��#�Jb@7@D�*�Â	Ϩ0�
9wd��Q�m�O
���>5�\Cպ����噐�0�'�����k�KT;Ð���-�EU��v��,���ń$@�VܦZ��$�QD%4F��YH��H&�G# ��i���"�gS Θ%���� n��"��?�K#��0]S"�&:'�{�`�	����Y���.A�?��3R��|��������vQv2P���U>�ǯ��k<�4�U'�̗�[���9������hMJ�`�SOO�������ysq�Xe\����uiq���T7�oM�y��ݏU+Y}�~��W��� ��΂AS%̚T"j�m>��Fb"�y}�]���FqϚY���{P���~��~�&������q��]H�'��#�C���8��8�+��@ٚ]��|�o���5,]��uBO�ӧk 8�w-H���p�'�^p���I�����_���a�/�c�%L{i��f���u({��?�LV�a�����j*kD�G|��~��
�v�@�F�9C���̫�TW��3��o�m���t�@���|��B; �w��?Mހ1�ԥY3,� ����!VicՐ����ğZG��=\5����^J=�)��D�I9�����W��XPz��\K+��xFyXNo�~��L��n�Y��2�Ž��* YPh.��s7��|
)#�[��=Q��\�ڋ��I�6������%\~mK���#�ߌ&�CQh>�߄[�K�q��{��O�(#2��1��{�|�DN�>1������Ǥ�G��q�:���x���@���ƾ������@�z�~�o&�uf�I�xFJ�����A�:̊s4����{ͣ��h\��
��L�'{�b���+����6���n�4�F�<1!�]�ڐ#������ � @yy��8L+�4x��{�H�������vNc%EA�l��}���UsBq�Mtn!M��-x�*�y^�d..K�OX
kft@��!�;�� �Dv��,k��]���)�=H������8��LE��9&�X3��+��d&jA��B��&���Y�1
 ��cb�]�4���煵��a������PZ�p�$��f��F�'o}rp.fuc�uK�����&3B��G��
���H��ʼ�� �`��� L����UU��U����̉������n��a�slW�R��G������8I�/�[�s~NWB���~-����p�%���b��eLTrB��2�]Y֫�d�o�ģ�+q�z��]�w�V�`r��4����(�����m�ղ��]XBXW�� �[I��G�Ē��ངH;�V�5Eǹ�PU��Ty�L� iLV�	����ε1B��Wy�=�S�J�1��`��G�Zk�5N�]�K����Ę��3�Aǅh<PD��#>g��X�����D��vD��A:�a?7z�K;���*�U˾�N�=��o|�T�dH$����٨��D[T�92>�tw]�_�AƦ���N�W���%���d��8P3^KQ g`YߐhUܛ���HW��S~�
���ttޘ�+��1�H��F&�̧�A8����T�=<;���g����m�.¬U��LE[��L'��*�J��5� �V�'����6❬���' �9;2��h�5�5$�c-㡝���sbAR����&/*Y�֋�Se~��^��p���ء��7�׻�s��Y�y�Dt�d�����=�f��r���n��ƣ��q֊A9j��d�3�⪍�ƟR���^��,�xk�73�;���x�ѧ��)H�|o_N��zpF����{5Os���؅�4C3�����V�2��Ս����N�?���+)��w����t�(���ˋ%G��2���
��w�	�������\�ƕ��:S�Fr:����/cu�,O��Z�]����bU�^��"qB���Ij~��cIb� !�L\����'��M��Q]<�#����vތ�]"b.����飣h���+�u���@�3�Se���@�\l1z�~��C�6|�SeM����G�8�ȣpR"�ɩ�4a�L��D� ̳G>��Z��q��� 6Ucp����^ _We�1i�Xl�?%��=YbS{\��-.b�-u1�{�WS��f R��/u	eV]&�t7w���^����+J��35q��s9ﾣ����t�9Dx|�zP%+wZ��"h����5SU�LpZ�����Є�~���С����'q�i(-�`�W��Ur��u�%���oZ��eJ������B���p�ܦV�̱P�Aœb4b�(����+Ė#�n}}T�������՛C,��p��� ���0�c/�ffp<��<��y�ԫ��펌��� �)���.	0C�@�v��H��'>�FN����u�C�N3�I�go�X�5�Ы+���c��9�j8���tdc�V�	;�c3��l',o)r�Gt5nRn�~�%5��HE*:�y!鷅"��޵��J�y�p�%W"�$5����;���Q,=��0��qwg�i@>����[�H������oU-�g�H�k���hZ���Ŋ��۸����پ�4��vV"i�m޴{-f�	o�2�ٺ�+n�����rX<��Ȗ�-o�^|�z�n;��<���V����������b��e��� '�Q�]w�N���Ǿ��#oN!y�@Q(��=�u}Q�G������r�������5�m����s���������v�m��W�����:?�֭�><n������al����BO�<O�zץ��e}�L82st�V �n�0B��X1�� ʹ�7&���Uj^��,����'�?Sa��E���/�p��g�w�˜��dd�\�qx)^��O����B���$
����3��V �n��ݱ �H~�·�7�>�������ߍ�{�FgDJ@ÍCX��^���N���$1?���#_L�ˏk�%!א�PMCˆ�m�#��z����h��y�NO�[)���@��n�nO���O�_؇�ؠ�_�)g�̈́�\��%�Ƭ����u�\p�c�'������.ӰƸfK�B������@`��5=%p�B��3���?��7P�2�!��'u8�w�:�5�Ȧ��m�1&F��gV�!�#>h��Mr�������☣pe�R�w9T��?/E9�����r�J�CM��YAc�')����{����L�����"��]�]m��3!��%��Cu'��aGk���H!�=�SP�q>_ycZz������t�i����7ٚ��m��JPC@Q��@����W���τ�dΈ?U�����c������@�֜,�T�K���2���"0�U���ѕV���$P�ׇ�X��f<�=
�j���W@	p:Ƒ�롇�/6J�ʵ՗�͇5_��2*o7���v4������l8�ɋ[f�Jy%@�N7��+)��^_�
n�@�H;�j� &�Q�C:\��,�^s�=��(:~^&h���9D-!�ξ��IASh���2'4���C����97��%vĖ��}_w�'F�{h��b����ڰ=9
�OS�?��4���6WM��r�;��2k������-��O��iDoC����G�,"f��` ���y��DR�������V��.e�-�r4���9(sl�n��4Fb�'�I�J�R,��g�ٍ;T�x�ܤ��YӜQ����oA���-�X��*�(h���կ���~t�:��ό�.��M�i{Lo{�+}�*��._=�+~ygZ�L �mzR�o��*g�әގ[i���=
����C]�^���Fo5!�ꦴt�-E5�t��-B����@I�F�^l�i���|: Y��`pŧ^&ʏ�T�_��l�D�$i�M��|�
�N���,5���-�ż�]m��B����}5���ޱz���F+���i�8H0Y�����ab��I�����$���/(���k ����dSJ6���N\�ܳ-9�5���m1���$FN&w����%/Z&�����s����x�ji�may~Q�9�3�+R����+9[�.wr�3���<�i*a{V*#�5���I��+b}�n�'�xPH�H���^cb��lm=�ُ�XT�3�^�XM6剻���̟��2)yV���i���GG�F��J�r�i^��e�y�l�u��b�e�(�%3�L��|�'����@��p�C�M&�bݨ�˾��h̥�a)��SĊk�O�'J��tƮ���	�:~:���L�%4�>U���T��-��m֕���\�VjVn��P���D�qI����ę_Ά) ���1���o/��k���am��|�����5�&@3U�ח3]�:K��!�*�~s�:ڒ�g�]���<}�_y�(��Gt>aR�] >;���w,2����|��Ȧ��Fף�Ꙫg���^�rǪ��\��<?m�2߁r�(N����"7�X5��ޤ_��j�G��X�*@�.�� ��w5�����Ӫ��8�t������Re��6	N�c�v�x�)V\Ұ*���Cw.޵^�x�fZc��~���3ܬ����A�z�6�*3�k5X�*ޙ���
��1�P"+@-������(y�x�^^����e$.E�l����L��}d=��"����P7i�;d�d��L�t2�G�|"�>���mi����N�4>��F�ð��KGq�p�K���Ȕ�g�є��5	<*��Ԗ��m3	[�N�Y杖��T�ۣ������9����jeY�w ������/�(�����Y��\����
�{��p'J��(�W@�����ߡ��
ͪ��|m���i�0h11ԥ�i��phA�*-�k�k���PO�5��GL��2w������*��=/>�H��W��Ձ�}ǖ��#�Nc=�����S��N�$*��0�Ա64�
��k6�}�vc9һ��Ub 6`M˚�EE?1����ׅ�ō;�Kp��>Y�&j�5����z�^��!�~rÊ���Px¤��@:'O��g��9R�����&M/�`>����6� #�nn�'_���i&����|C��� O �8	1\e�x�⧋wA 
�L��v�"u�v�ͱ���?/ǡ��Q��sA������቟�h�L��!�πy>��
�.����qNo��RǗP������;du5�58y
�U@�l��^�=�Q�����k���`�҇h�z��ɔ��*-�o��o�C���V2ߵ�l;sI����e��0�|�$bG���pYEIr�I-�X���0ȦiX/������&g��+���F�� ���Cq��y[�3���du@Z�?�"�b`?R,��C*�U��'b��z�W��؀�&�@,]ĝ�W������=2�Z��Q�!�?kӫ��:�?��4���Y��\�Ib�	:C���E�O�u����]} �#���䏟P�>~���N�<���ݰc�����1'j+���*.�A�(�h��=��I�,�)�CT�981tG�~������#�d
�0L
"o��K�{�����]���	��MG�����/	^ˁnI�B����,�z=L@��TN�D���ᎇ���_�.z�4�����Qc�����!��C�lܙ}]�w�&�.@�\��?4��?3Mr�޵���,Ϊ�fz����z����C��A̤[�t��!B��a�FjRV.�2$��md��N�����,�u���b�M��������Rz���>��l:Oe6��2����)�&�GC���@[�4I�^�G�ID�5|N�A۟�4�e͘-|]b���f�Y�joY��w���WS�8�tuY�9�E;Pxv�ڝd�����I�5�3�ߠ�P�n�V��+���t��ι�KY]}��h�\���o����&ع��K�p1��,�0��*y�C��M���o���N��&:3(T�.�X��PH�v��MJ&M����U~!�޷�ǟ [�U�0b(�E5Y�-	�����2�=�7R�ȭ+�V�ם�/%��<�²,O_CQ�]��={P�q0"�tϗ�x�ރlI
"6��y��#a�)E3W�3*0��C9�A��P�c��D����c�P��h���=l��'1�J���w�k"H�S���9�e��
L��51�������CT��mt�h�_w���V�J=�̄���X+$�'�"U5�:�E|]����̪_	Z�1R�}P�����L���Q���rg�E[����D=|���_�M��B�]3oR��*�@ɞ
��>���g�.[����	��].H��0����B�C\�K��Nmk��_��fF���zS"O|�Q}3���Bq�OɂZ���L��R�f���d��c"��n����lf���صR7�mk����R���z���Z�4;�%j�����Ď�\�4��$�]�[%`��!�d2���f�DzA��@�i0U5Q����x�0����p���{�-�� :~T�γ����o��B+�j��7Z�ͣ�K��vn/�4��!�h0�㍌N�>F�Sk���e0��(���t
8@���͞d�
�\F�-�!���k�>��:�����imשY�aw9��M^�f'޼�O��OsK�tF��W���T݂˞{��=8�v��7�޺��-����J���=g��Q��ðd�DS�2�lr���b� �t��'hn�?�̐�6����oà%BJ\��w��N,��+�t88}M?��ac��F|:�N��_~D2�Q���^+Q �T��6>֮��J봎�L(ځ���r�o�Ҕ��r��ȝ�8���W�za)$��]�?� �Q�v͇�9zI�m��A>�b[=���{ltG�`�z�p���])s���tn�UJ���EbVه�D�}���ϛs^��7�7x�>����rB-��/�Q�܀�����vuO�_��?�d3*[�S �u�v�Z����Ŭ������ ]d���ۀ�2�k�"}�>=�P��åq;��5p�,7����3b���-}F���vA��T��, G�*��vo�˳������7���_\�[���b&�Q�ǁV�R��8b�oP���"@����^˲۟ݷ<�I`���@Z=U�kɛvW�<��}�DpqU-���2lg�T�qٌ�{bX�G1�7q��y������	 �H��:�5�s���OϹ�N���Q��0��ɗ3��{�鹟�v��|���BWL�/2;E�?�pdnMn��N�k�V��*Ŧ zO�3�;�z���UQ��}FR�� }a5
�Uy�]��qf�'s���Y������\�'���J��M��8x� �.�G��o�n{�(��A���������L�*�m��7.��x	��!�2�Y��^�^���J��-���u:KW�0�p��e�`;��q�v