��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&�
TB�(+�
mQCJXk�ɒ���S�H��U�(�c�H�u���\��֔�PW3�-Ƌ�!���A{���X:��fu��6}�#�����X��/IPz3���y�.w�>u��6�C�
8�x��^.Tq����rF덷�a2vBv���!.d83�,��W	r�����w�NS�kYM����l�L��}�9	k��<�>R�a^e�&�:�*�˻C��ᮮ��n���,��B��m�Ki�1������+�9�D_A�=�1�C�Ͷ:�8�:?����#�M�(�<V]lU����%z��FoTN~�~!_�`%��V^�}�����u��q"��*˫�UHm �uz�Ә����bKr�]�6`"!j�Mr�����Ī:]9�X�P�UJ�����(�%���k��!�������YSJ�s�ߍ�k�J{�=�Z�֐�L�"7�P�� bL^[�J�����+#_9�S�j�QF��8��Cqe�b�F�uVtjC�N�� �K�AC1�M��/R�mψ���3�e�GC���J���Um����(�i���Q�gcW��e� �1��Յ�y)��$+ ?�'�'���CZ��	4�2N�v�@�$�䯕{��d�QP�'A�I��}��{�_��D��+�jɪR&��>�#Q)�5�b?�,�f|��__��
�o�x$s��)�l�w���gA�S��F�X̖�B �Z��e�,̶q���b��șdM�E���V����`����h�~�:���a� �dK��&xo��@'5 S� ��������h�#��1ί��y5��9��xG�$|�m:S6iY)��3iE�^��4�.AɯH�g�ak�PV�~�t�ѐ<������:OC}au	��&z����<�|3o
�(��s�	��{A��o��s[�-,8g�:�ڿo,���5���X_�vWof�,47��y\*W؆�LL1��mJ���%��X�)Q4���fA�ʵ�|)Q=e�L�#|��9$��6^;�N�=�d~��: 7�n�'���������`:[\�H<J>-G���Y:�;�Mri}dq�5��/�Ḝ�T`��^���"?��{�8���%��$��=�f�fV� !����X��
˭gG*jBMb	�������z�f��o������$dP�sL�ڐxn�ڶ�o��.��a�N���|�dҠ����L��<�bnU"I������4o�	�^H�ԯYFDYH�W"��A������B�W��6Ŏ� ���.K��.6��%*Z�([��0�

I-�-��tg)C=D�K��5�Gd_Z�B�=zN��A�J�=7w2�}	h�͐�Gk�%eh���	)Q�$�Xw�h�S���ǌN�61����ó��3�Z����>�clr�O�*����
�j>T?���LB�Y^h���;WMWӀ̈�n��]�piN ��q[�J���z�Y�}CoG62"�x��0`�\8�"�ӫ�cmN��#U^��;�S���!I�aÛ���^̙�v��'
�1��}�{�3A�
�������1��3��{��J���k.'J�*jP����$��'�[sQ��3�1l���R1��v}�F���U!�js�#f]�1���Ja۷s��̊M-�@i�_�^���]T1@�J�fҬs�G��nZ���\�
r� ��؀ߺ�kk�^�����UE�NM��m��yL�=����-��"/x����n*3� �@7Y���b�N�X��ܱ+Cqg��n�v7]���18�듉��P?��t��W���	qJ�}�=��+��Ia,��r�^�]���m�y��;/H��{�"x�s��͠������6\�J�I�D���l�k\7�.fBÕ{&.��
�JB�7f��-��Y~��,+�i-��~����&�~��G�Y��:�O�5���D�N%����{�n�n5��^�	��>w���I������:r!-Ϝ���5+G��b��0���[�^{A0��h��;��&�ਠ+Z�0s���{���Hva�oI=��7��l�D�X�	�^�%s��[�t!�Z�f�(�>��,����ܾx����H��m��>a�� �U�F��U�K!�>��^1L1\@ջWE�nc�Z�I��j�<�8�����?*�����v�'��:�����.<�HV_�S���*��_+S�H�/
��])e�)�Ro y�P�2Æ��Cq���(��1?�DC�Z�3q񐝵��XNϙ�L���=�j���M��P�Bg�|�9��8�9W�/{. �c�-%I��ORG�</Hvh�� �;K���/	���v�{d�wC=t�vo}�D��dIG�~���iل�� #�d�Е�����_:�g,1�	Ϛ�����u���9��K,���\���Մ#�?φ&��W�͌^������2��Q;�䠴x�اJ�u��CU�����:��8֤@�^�O��(X��p0\�j�0�چͽ=o�G���<a����Ui
�|���+˒��y��G�Bx�����oa��v�>q:D��Q�)ˤ�(Z��{���y=�j�;;�R2A"��}E9��hS��S(&G�AM�؅N�^��5/��ɮь`��n�����`q�M�T6��L�VUR8��ʽ?/�-
�}mv�^�����g�	����i�ϳ��JmTL��F�e��m�c-�
�&������sr�WܓҘ�e����?>~*r?�R�LG&+lW�&�N���i
C�p��y`G�om�����M4�G��	��}��UL�I�/I捈Ĉxz0�%a��xm�^|0�����G���ΣP�ͤ���.w��ڶ�;{Y�MY+L=E��.�7L�㣨��W!ek�JO�u@hR!�I�ƁR�Y�z���Ρ���d��\�^�S�:�6�6����N|���rF�o�9s���?��d�bc��hV�JO�IoS�7����J�Q��]��wJ'�S~���|T�xȨ"��-�l��U�3 4�>��k8=x��

�+�N,�+g�9>*8I��Lr-�"��!�Jv&	��	�@$��48Qj�k_���qϩ>ͽA9�R����k�@�i�~�;����H��1��4�mktp���� K�L:Z�F��`�Ew��>8�(��Z������mn�[�m�{�י�O���;.Pߘl-V<
e�r#�7��AI�;�>����.�ӑ��n��K��:j�l��z`�-�M�O�X-��R�$���>J�em@�M���?�+H�#�5�����rPۖ&�i������� ��K���*�1�p �P��ay#�+t�ʔ��~��d�~��v�<H��h�e#�L'������$���c�z�S���5#F�u9תِ�o���8�i�~4�
T�fV��;���?��E �����)�"�*���O�s��!�"]hoS���!�uz��b���F�$�^��c��}1��A��(w��j2����[I��7Nw����5L���q����Ͽng�\8��dJG�� �<5�E���*N[����ߩq>E4�F61K6!�R��.�U��6�?"ܝ�^NІ��(��0*���^}.�Gg2��ԿC�����'H*���2�|���4|�����쇚�е'�S�aZ&_���-T>c�6�t>�`^�r�$>Q������_b�����0��h7��shI<EJL)�AS��a��@fR]t�3�g}S5�,BCf��W�8��[.�c�ZX������a
F������E��q�����޺<�'�"����CY�0G#.�9%�(�%��J?��;��OG��z�F�H�3��\��ꘫV.��� �k;�$��u�p�����������_�_Q��C��Ӝ|:���\�k�*d����<��y����Xa��B,�*\Am�$�;,�=�T�|�U�V\���.�r*����"k�Pע�5��XQ�?<�^0��� �VIn$`��IT׍��V���[� qO|�sa��[��a:��d#�1雖�n��&�W��+��Q��*+�А	��㍧��nSr�ׁI��A �x���<V���~��T��t/����
0��48@��̦6�f;��VN\�x;CD��8.�����շG���aИ�Y�ed�����ew,�p?Q~Fځ�)l�X�k����w�e3����v�� EjS�H�-�d~kAu��N&�W�����Т�i�p�]�)?��/�"�苳
!p����-��V)���$��[nS��9�:tV���"մt;�+�j3�5�AԚ��i�0,l/A������\������0�9�2P�vې	 �!���A�kPBP��[0�����?����U�X':�QΘ-n=�L�%>w�5�(�(��߼��:?{I�AO~Z�e��ǿ�)+��%L�v �8J��Rs7��a�{0���T7cp �F�e Zh��8B�f�*�~�����e�͇��V!x���J�ؙ��rUU����1����M�x����zz����܆�+�Ԣ��9�;I��md�Jd��?�_�P��h��.q�.�
5�c�|T�F;b�K�@����v�j��I�_q)������ǟ���0\�.���(V��ǇK���[R7�?�� ��E��]ԤN���r������vR-�Y4@�>��T �s/��og����0���?̔�-7 װ�St�h���ԍNu�]&� ��-kS����x���sE��vz9��/�e�(�]ҼR�R����\zǰ=gi�??D��xIuX%3����GVeW��ZG�I����2eF�K�p����݃�I]c���	RƘ�|ִ+�]�+w_D�>�3Tz��\"1?s��r#��N��E���n��Üp�������}[n��9�w�.^���f�/6h��E"3����f�T������*]{؟����7)���p!9�E����"0��>�a�L����2�3F�+HG1�Ƣ�}���*�w�W�W&W���c��4��Y�F�ڒe%�����On�S,H����Z�ԵF5m����,)V-u���:N5�2�݆`�B�dA��-�̋��P�}���=�,�:��e�!��kv
r�gs�:��QT�g���6����0���N
S�e���ĭ�Uv�b��'I:S�f|��=�9��Vsm0�xf兡!,�:���ɢ$��W�n�����w� ���d�=
���*�0��/B�>vyJ�7^�\���x���� OM���2�dۥB0؍\t/��y��A�;���g
-���g~���P�#@����.F�i��!_ߝ�켵�a�.۝׸�&���H�u V�
�D�k�&�������t���K��Cy4E�ş���Yj��HBR�|X�R�PA(�c������u�_Q-v�k���p��-�g�4
d��b����,eF��%����%:��v,��ʙ�KӔ���v�u|����=�Y*t0�[�1�] ^N���rp;���������L9g��4n���N�^\��Q��^�7ؒ�.B�y5�h!(p�0Ro"TL�[�'���[%�_��� rA�����~PI����:	^����?T�h��E��@�ē$Z��B�+V7�����b�/�KUz��i��_��4��#�������4��ۋz��n�'�X�|<��;U47xK兓�v�N���A��#jꔰs��|��
Q�) J��Q2��XC٥�q�wJeߋ��%��72P��#�������{ ��ݷo�;w�>��7������Q7�]V3��WUiơ��|R�����r�.�r�1�@�k{P�R���_�v�:��G�pq9[�e��+����.'�A�f�į�+�@b?�c=g���%�=��V��2����{Ĭ��e��Z�;�$c�,�]�J��|5�<EAu��� �2�4�e+���n�M4X��%�? �"·��!_���)U�h݅�N��L��)熓��D!��K����.�w?M� /��u��oLa�⨘T�H���#�l��KŽ��h>�b����������ȌD+���j�� �`�oi�j�h�y\�}�>2V����������a��1 {i��?5[<��7���d�)�����à@�b쩓5w.K���up�'�	�" \�Z�⺅���c���wV�C-{��;�b�Tupѹ���]`��t
h,pCGI�i�ʔsE&d')Z���Z�	\�ٙ1C��e��kE��q�w�!��f�mz�U.������28��N$��Ur᣽�sK��c�E=��]z�-�P&*�&��U�&��gi��ߪf;�=P�X�Ӎ���0��͢������(]���}���4~AM,y�ѫ^⸂q����T#CI����O�DƇX�>�LJM&E�/z�5�.ɜ�!��*��2H�����"d�z��4�q�ADiH~��������fP/����!�˛>���Ҽ�2"]��$��}���D5�$W������$	}�B�c׌�x^u-#,���n�S��`���٪m�}+�c�@6�Vlj�漖dƛ{�):PV����r�[����y��s���Z,�k'��"�u0�P��/t�̡�4�0(C�ӝ]k|�v�|�:Q�L�pX<�k��ET��dۥBM�5�����Tys�8�>��M)Оџ��<pN��n�!���
E;�-�ջ����`��l -Tg�S��ߣ/k�����Q>돾WR�7���`��L�6KVv�������_�f����p��5#BT>��+>7���\6�� f/��]g���bq�2���As��=9�o>䠞;��s�~,
U��H��a�i0o�:N�ɼ~���.�P#����S��_��Z;m��Ǜ>��'��Z�+O�mf���H�t� _0z��>�}�I�J�H}뙱(����s��56�e��W���(�nz���fr۴��X�!�aSv�;i
R��qī��>��z�x����,�e��KО
?U͒�QP&�QÛ�:��%@���g	,�{N�^f��8L�`��������~�(X�mZ�e�~w�q��Af!�H�".������JS��
� �BA���N�U�~��X!�L��`͇��4v���_*"ܺ��O!�{P��S�|��D�?�Ef�Wtd����-��5〡�O��O��Hwdr�}�d��u�p�7��ȣ�W�|*��:�̛'�B��-���qp��Rm��[���Ò��>)�I@��c$RW7��%uDn�4*�\�>)�q,���d�s`�	�*�D�kF`�������=�՘�C�s��xY���2A���K#��_��gi�����H�+y�;��}q�P������TV�Su[�a�z�"e1�K�z�\tݳE!��"�{���Ɗ�����I'����e���mD�O/1P��%|�^��&	)�]��ϙ��\OTQ���d�aX�rq��@�Yv��ۗ$�A�ϝ�d��c.r�z/�U� �P�o?W~���	}uwR����v\�a���ځ�i���6�AF� �r��~�Rh�e�eS�&��R��ὠxm�Z]��KS���4(��:��B7�ǚI΀|�x]l�b� �s�%U*�-�&�׺��qpy����+�h'm�;�i�G2�&��G!���(��bS�4�DAǖ�Η�XX�1)8��Tȯ����躒�/Ц��o>���j�Aȸg� ��T���A���(�f�u�Y�h�-!%��PWS�*^2�\EW�eXu_�&Y��\ �!m�V�)H[�P8͜��qS=F�z�V�n�Mi0��y������73�f����@��N�UKQ8N�]t��F��\kG'�j1�AT�j�9���oCf�t3�Q\���L�	�Q|5���Jb�%M-��@� ��#�fc�� 4+D+����׹�u�����teiڣO�G����ćz��l$Q֏��D�t5�y϶��1���f#J]LL`Z�Q��(,(��6D��I'�^E�̯Ǽ��y+󍇰����l4K�V�!y�|���2،r����2tYΟ��FP�	2��b� ��E�ft;�p�R�Ut�v�	ƌ���U�7-i�h#ߎ�3m�����W%_,h̷���!W`S�����lx���ƿ�J��<:��>K�ס������������zL�g��Q�-YqEa�����	X�����pWw[�>L��� �/ǭꘌ�4�Y��}���َ?�>ɕ1��/�C����rH�dS�-Z�g��ܴ�ڥ���F�"7	�ҍB;���S�_q�/����M8	]_ٜ{��B���8�V���4�ѫ��DցGꊀ�.( �OE��o����'r� [����(ň41!ǥ\��)��<)���cH����X!��,�Fr?E]��f�QZ�?��=�:~,�h6��zr�E�ZL4\���h�G�^,|K�09!ڇ.�`(,�n�'�=6�'���Y#�ֽ�����ⲵ�miH�K0-V!����(^��k�z��ph�>T��ҹ�c�@M��g�Q�eR��|Ź���U0!���3c�5���q�����D����jtYb[�RDe��91E���F!�1Od��d'Mϋ����<е=C�du���8�`��/`%U�j�G+��V�
5����u��_�3R#��Ȯ�O�ε,�dvo
aW5^BaB�oů�}L�>�>4��� i�I�����⁊�/?g�[	��7T'ѣ���A���wM�Gu����'���C�E���kMd�G��fە�����_oI	=H�N5��\��@��K��-�?V%;�L�)��Y[�=��<��+��ܣ�/�S<V�X���n��ϧ��։�8f��j��KQ��al�sD9	)W��@��� �����|:�P>�	[2�������[p �q3Š�Ym2_�yh� ��G��N�'���Q�����;ӱf�sƼy޴�h�D���s�:V�	�.���F��.`�8�뇟O�HWF����n�t9?�[�-*^b+���[�ړ*��T���iVѐ���VI:��ʙ(:K��գ�j��`\����T�� [�>Ͼk�����QnF�ww ��]_I�4�C�*�:r:�.�5L�V��6_/����=>��1��.��Xw�9a{����U�')��.���7��a�c�e9�_��ʱ��㨛u�Ŝ+Y��\ˬҾ(6J��� ��^ly�'�СC��x�Z1�^�9ك���k�`�0���{l�N��/��C�-��h��?^�v*��x6���֮�]��6>���::�Rm�ay��}ђj+?
.����@��UԵm��38��>��������u�:A���Z���0Kw;����X,z���"���Ռk�l�����V�E��F�F��@�`��&�r�g�u%�s� i�[���Xg�
.^�r������u�tj"<��*z�����^| �� ��������$ì1?p$��1NǥH����ȣ��T���\���j�+��7�S�<3
*�3:m7�`y5�C�����N�m�W�OnQAx2�Z�P�~�G/��y(�a +��*���E�b��B?���}x���S
l�ֳS0����$�l����Rls�u�Sǆ9ʖr����8?S���3:�F�����_q��aSkb��>9tUPJ
D�x��χ�.nni��G1��1G�oQ~Q�B��U4�V�Uӈ�?]/ַ8�KL���n��P�x5ٹ�����&�nӟ�]�l��æR��6sT/� ̨�<m����{CA>b�z͎z�8���R����I�8N����f:_���^�W��";�)����
��(�2$2�#�nsP��b�>��;H;F�o)�������:�J�^5�߁���/喑gy�g���0�����'ʄxN�!ڣ��xM�{3!0��jhS�sx��b��s�D�LsZ�~��I>?���A�0�Ϝ��-J�L�Ʉ?͟/X��k�"Ä�.֓, ���w��L7����3�8aL��Ց��<����A0�1�t~��,Iʰ�<�n�X�|3�U'���cD�QgOc���F|�3���h���?<��+�nP�B���4�����C4�K������sǿ��[�%*�D�-�O�s�H��Y)? �nٗa>y�]Lu.(ܚ&�mc����n�፟�,y�m^e�E��4�`�֐RF=�*îe���u�����DY�A�A�}p���Y�����z�@sS��\�ѡ�d����j��G0[A�o-6یиi�kg쯬���ň�&��w5�H�[���>��� �����9i_Is�5C#Y~�ڪ>[j��9$�*�r��ӡ�VQա�^TL�A̼T$����׊\wf
i�6�;�a��2b�7���#h���pM��y�G8�d��@���j�x��]�<�b=t�N�
*����8�P��yK����T�r ��bZ�6�����ƥ$�>��uS�k�D$9�C�T+���x�k/�G� N�Ѷ�]��#��p|��â(��v��Jm��ގ��芕����އ]���J`�X�k�����n	a��·k=� �l���!IQu�4Q��cA�\� qe�?��J�Z�����u'R݈"J��2�-$	�w�a�0 ��(�� +/}e�����y�+����QF�R�x<'k�0�\W�0�ϋ�Fi�|j+$�ӏ0;z`�U4��!z��яu����#�������A�o@/�_�bHX��h��u��f�5i˂���W����`b���&����"0��3�c/���+�N��/��{�}����¶��Ѵl����#�jcQ8ʕp���+'~ϒVGTZ~�L7�����8DR�<(-
1����;r�b�I7��m[�=;g����)�d�!Z����+jQ�	����K4$�٠���+J����W�7�}T̑"��(GCb	�����o�GR����L?��]�#�U�*��=�"�=AV1��@����W�T��5��F63�q�ΰvS�("��tCߧ��Y&�0�欋~��o�H��𡎼+��F�vX{�M}�2�yPF9���jv�>��ؐ���K�ʀ!������n�K� �����r��J��f���N�0�60�i�I���i�rQ~�������P#J��0�؈A��1	*[�"5�Q|]�E2�$g��g��0 ��&�����T����Ґ?���h�<�\w�~�U��TCv*0-p\`m��]�^�	3�����:��U������+���:P[4�¤�~������<��0����h\�]�iPo�i�X��2����R^B��"qڈ��du�{�7:3�������%O0�����h���_���Z��cE_Q'P5���ȝ�{���[� ����]#���Yw~2l�2����S���Y�O����4����i�;����0#2D�.j�Ì�J��ѵ_]����6L��<\�{Ոd)�LL��$���W����|m���>�& 7�u�\���E��Y�!}�Hi�{�o�������T��}33s���V�y�:+Q�$�5
�@)�����}X=��0b95V��x�� _�6�W0wm1%�~h�L���,���|��b�Y�=�vj��&kev�ҔfvJH�P���P
�`���__7����U�(;MGc4a-I��Y"*ӫ#���֧���:�rS���-Ttm�̅`G��C���4��C˷]Ә�N��R�!�4���=����$�A�?阾q��� �6PIt��o�|s���o��/�*9i��4��!ہ3Q!otӷ_\�<�W�T��g|%g��� ��h��鞝���__?�m?���q6|$�Q���H�w�����΂��N0���v.��/Ĩ��G#zk �`]1��������{�����ꦰm{~��
c��!"E�g:4\sc�����R�m~��@z�\��[\W]F�TCf�cWE��9�	=��~ؖ���[�>bi��+�j����8P
���9�ߟ�i����U��k?�9�Xo������/FdF\���Q���F	�e	��e$ �I��i�VB��H%�v���QJ�� ��Ľ6�߂�IH��*ˎ2ɯt��NM��˵9�f���mz-�M�� �GP>��XRA+�����LgH�7]�xoAl��*���<4D���F��h��I�nJ�.�J����^� �>b�T�>�R�K6��ap՘ ���\&A��tlBHk^�-,�i�y���Fl�����v.#���k�!1���&�Sb��k����u6��iK;�2Os-^-�즏&(�R�㰲�e����[����Lz�t�)���_�ڡ���}��_�ݵ��Eo�`���l��4���2�Ҍf��Dj�]�n:�yЊ��q�W:π��1� �٬^���"���([�44��d����b�� ��'/?K�`M0��G��4�: �6y�54=�*^5팁��fy�;�J�_�R�I���m��s�j;"|�6�����V1˛|�~�%㎰��������ke�$ .��<)�ս1���|+��?�`[��K��Ώc}�-��@����+֞��sA����8Q_H���1%?��e@�.0�= Zr:IP��h{4hM��F�I��v��@x����շ:|�@�6�I7~�Vw���rG�,��.l.O ���kQ�������6�J����F�^��H��?��(ZFqYf}R����V���b.߸�J�ߔ+�C��]�`�[�]	�\D8�s�}��u?
5����Q
u�?q�C3��0�E��gPZ'7T��3��΂rV>f>�eaE7!̊�L,�()�m�DRI��j@7��pY�Q��\���:�H<R�)���k����8�-�Y��_�4���3�V��0�T�!�7�\З���X�]��>�V�6��������]��H��0�ME.C43X�ʧ V)Zd91�dr�8�˨�T ,�������~�'�Uپ�����8a�j��� ��&ձ���e��w���ϵ2IA�	ӣܒ�6T�.�tV#��z���Ι}T��4�k��tV ��_���B�Jl�����.������)���g���׫}8ܔ3�&��a�H���p�E+�Ui���g����Ft�=�S���Au�j�5���A��H�L,���\��'7j���w=w[�:�L^3�`�\ǛY� �r��;���Tٯ�w�{^�r�2 uHMs��A��H�i�����E#-9����
K�u澹&�����c�DH������EV�VW
�y\���9d©@oʁ�e�<�*�s��q8W'�:Ⰿ7��Q��Pn6�~M��]��C�����}O�c%�$Es��I*B58-�?�u�tU���S�/�?�).ͤ%����Bي��� ��wkQ�:o���KśC�ʴ�t@F�}����4y���v_�����&x<��/�^wf�k΍Iא���v���$MX��l�;��ه�M��7�}F˥��)�1��c������A�>K����4 ��-(��0i�g�0�g�B�:�״�� �K[=��ࠃ�(yl"��x���)�F����쁡���{��^VN��u���&�ᾡ}�6��Dm�X��ّ,7�ѵ��鲾�.��������CQ6�+�����]��9�;��Anrs?��m@H�"�Hy�����X8P�nR���N�І�t��%�n�4��vs�F�B��}�����Ţ�G�i�S@-���_J��<E�z'�	��H��&�w�L�J��S�0*��bQU�1�x��!%�d9]�f�B��-�ơ����C��r���"��Q:-�~.�}K�jЁyQ�.>��SrFJGc��`[��"�� �&��2�T�&V��A���C������?�%#��2-x7�g	�6�G�����)ª�H,x(E�S�ӤS��K���5藚�T�E'��]��Y7����k����̜a�C.��a6|Ŗ�V�b���/p�8��Kf��V�C}�#t�p���m�ES��<� 1��"a{� <<￦���!��$����DT`Yb/��h�C��e!��Q�]Q�u0o��H4Rm*�7��uK~K8?!�ɂ��w�M��lO�n�W�[���%�S��x�^K�n��x�.
�ci}F1���B��j�h��'&#G�Z�+��(��]�;3	�$m ��^��v�O�9�>eD�8߉hf�uJVA��#�܉���x�Kk�i���3�.���8IM��旊�W�"/N(ͱ��"+o�0���Ikg X岤5��a����J%�h�^�t�����u��I��b �T��݄�腒��VC�PZ�S1L�������s�5չj�Am��YT��n�	��Ү���B�Z�E�8"e?{��|쪨CLBb$徤	���-�X�2�ak~�� ���-��n�$��|����qŏ��k'#x N��~$?>��]����KB����M��1)#��p�D��Ė�� m�(AKs\��ǯ��_h�.$c2LN���^B�<f�.��ʓ�>�e�#���!��1�@���;q�����wB��+�c�V�)������7������$V�n�'L^���NA �Ft�w�n8��j�AМw<�~uG�?G��j���|�r�k��{ �!�����N<9�0�gh�ʟ1�nX_aQ@;ɸnف~dW��+�_r|ۢ8�����,��x4���ل{���IipU�6��$6"��zv��{��-�@��=�&AH�	�0�"�¼�}%z?.�?eMb<��j`�h[��z�ҰW���w�]2BE��⌇�e��J��j��M�~n��S���6�^�=���D)2�ϊȁ�K*n���a�?I�E.�sM�<�u��'D��I�br
{�T�;btQ���ʑ1��x�4~�MP��}Z|�3�5���흔`�"��ӿ)]���>Ja�d��?��S�MC(P���'	k��rځW�����)L�ϝ��\_83�|���Sjb/��3Πp�W���!�AU(q��)��d������i���,~�*�Yc:�~�����ɿ6#P53�G�ߦ��!�mS�N���6-��(*Ͽ{��9+���%�JCh��oD�D�U�"�5<mEtmRLV��M�rwVcU5\
�Z��N��N��K�Vq���XB�+n9x��%��O��dȷAK3/JE:�h�|��c����K���.i�Q���Y�=�|>��N'6��������r�+	�s�S�N���{�*�q��U�,Tb�q�*���j,�SzZ=��Y~�/��Y�x{�i�d$��7�cY�m�Xf%<�� ���g��+�n�o)-����E�ʥ�E�L����H��`�rxڑ��_��h��~�ϟB�)��*��X�5��U���1�k5P�
Q�£�;Տ��u���C�#F�����?�g��1�|x$,v���pq���Xw�λS��m[�#�^?���c��k�? �M����2RE��1uq�au*[
�����$4�W�p�D�PjQ�n"�n��>v S	BJ}X��9�^�����m�O��Cm�7챶!�%���c\@WhW������"��v��dlۆt���宮O����ɭ;g�헌��N�9x�\u0��}�"��H�SʜHzq<Z��c��]��!�!+2A��'a�=JJU�M�f�*�N��)fblm���)��M�������È��o��_�ww9��������X�˷;i��G~-�g�:m%IX�?���9���S�����s����Ѫm>{��3�a��d%�S�����®'����~�h�Ş��O���vs���D[�����q��?��.�V�,��~󨒁W)Z��&NS�9�	I�ԝ��'��itH�������cΫѧ~�b��
����K�xqI����%�&&���-����3&A���Ӂ]����E(����,��E��O�s߃�5�R����mЊI��3CF{���)L�ga����,AY�2�%��J �V���&^F�S* ���a�FL1ݕ�A�O�=���̫��7̶eO�e�J���2v����=��Hmؿ����!���/�Y�9R�z�lF�n���n�;|,:%(Ѹ��~ �� ��a��e�Ʉ����$���B@�	��[Z���[���`��h�ix�����s���3��殙ұ�b3�'�] �����]���xݘ��%�jud���ܑ��}�"PB	��R�2��pXƿ�W,�{-z ��+��������޽�,�Z��|T�;���x)��XA�����	�O��̳L����[T�o�I	8�?٦*$ؔP��L�L;�(��@�zػ��ݮ�BCJ�tƩ�$�iժ�Y>�V$C�j�Y��՘	��I��&�L��k�u��Dlw�f�("]wk��r�� �H�q�Z�7\�>��7��4�w1iW��N@(��+Pζ�[x�r���OL���+Ǵ�3kr-A�@M�:w���f�a��p��x��\\��'U�Hrw����(�`�[�l�o]Р :��?6�s�+FAKm�bD��8q����6 ���\'FW;ܘ��hej䜥 �R��͂bS���n/j!o�#�~SZ9��?��Qc�k��T��W6�kmm��Gsh�~������}ے?ݭ#�>�WάϞ&d��|Xj�I5�-���Un��z+��F�n��j$]���. ���P�Ii�Ͱ8������Ԭ0#�����c����%}��m�^�����̀�����0J�������1�X�:Y�8�ͬ�l
� 'oJ��C�V�q�^���P*]��m��M��v�Q^��	z�:h����� �B_�x��Y����4���]br�¿ԫ�=ֆ�ANl�=$��y���yQ
�I�b�;ܾ���y&���#P�y~�2g5�;��� a�X����`bX���,� �z��QY&�u7�wƖ�7[��-�/�B6,�rGA�Z�����7�qo��uڛJ��'W��<g���1�Ӡ� �յ�)N�L�U��z� B�l�pXw�(���� 9���P��'N&m��~H��)��RLF
WM�r��S�ͮ�7�5E�#�O�rk����@�E�wM�mGM+���/q4���m�Š���t����}Q�aw���{$})|5O�p�$/�Y�c��9�t�xe�|菦�e2�e# �� ��^R����#&�h��`��A��!���:�O��_����dxɚ�|M%���i1�QvT�<.S݋=�F�~f/�B�SpJ{�_���VG��v��7�����ɿAJ˕��L�ԧ�/L�6U��X�`�JγJ�H���%	�d�w�e���V�E��8(4�>���r��^��/J�oz���!�"�5��&��X.Tߴ�qE�b�=H'=,a��b��Xi�`
aeǑ#�2-38a�s�8��"4�-Õ��cbS{}Ԉ���DPF�VfX99zz\��n#� ;��!�y�3+m�;�[83[ɾ�f�OK��c�i�ò�"L��)l#ɔO���ø_�zY��Wq�~׭���N�`��6�nR#�8�3��--f�RZPh�X1��1�x;hV �U�QH:���s[[O
���N�=kr7�BsxA6����F9���]XQYo��#���/�F>g���IB��Sw
;&�<����� 3�}N}����;�Q���Y:����}�5�Q��%�����4�#%g�z�&����N��S��D�}ќ����E8���� dCK�n��Lg�z�r|H.�i���/$�+�"��6��	�QF�ċ!����_e,E|gB�JQ��~�{����^R�V����XLc�K�w2�pB��/	�|�V�e��q�����o���d�W�ܠ4��#0E����ӈ�H����Ud�4QU M)(A_�P ?�������:��m���eX��c ��#����Q�S�c�G���]�_a��%o�I������`�����^T���5q�G�Y<�;�����-��g��H�n�
6��I��yYqyzgf��>Ԕ[`�/M/G&�p3���h����d��G�Qw�v֔
�?�DQG���ټ�՜��֥�-����C�p����x߽i��$�JP��BB��h�P�x��ń�z����0�q�R¿��}�f�9�U�䦚G����%r��s�3�^^�CM�5r
��fUn���!�!����Ly�ó�M�2Z�h/yL�h�-�G��F(�˖�ߋ:�z��G�*@�����\-k�rAI�,�$�<�J��i	E��ι#nA���s�-@;�/����)�.(�TM݅@j���\�d�p�z y��\\%�O�q�)��\8[ЯHE�o\�;&��Ö�zءp-"Ļ:���N�%�%�R��9��O���=s����B�̆Rm}�]�Hr-��ȥ�s�y��Iފ��]��3�^I��ME.�-�5�:mZ��{z!,[��Q{��t]��[����u�u�V�Gh��O����jZ�j�����O��.�w$�@��>ݵ�p�&���5���Z��Zޑ�ߺ�հ����b����{K�`ٝ��T��U�aق�[���Rt��Rg�Ҭ	��6�a%%�� �͜0n��X&�SU�L �Mo gZ+�#�H�rkͳT���F�O���ޠ�˨>f�E�*��N;�k�:�}i�,�DR� �����0�o�&WY���n�P/%���2��F���w���(��y/W#����b٨�+Zc2C���|�=��u�M������C���ۑ�ϒ�Qhr��
�E�RŦv�����S` ��Z�H�yXf��ʯ1���?����Ԁ�c�,�=-���u���22���WdLy�ݡ�l���*���QG���˾�Kt�0�J_�)+�yAW�Lj5Hպ.���T�)�v����|*���h�D�kef)��@���>�,$z�v��B�ݙ��_'o�CG	�Q�7X���?J��'�92:V&��Mͤ�|�b�u�V�G=t}��Y��7ɠP�����kA9C�6�H���)}�f���4�:J�\>��wE��my��xvK�CAҁ#W\�#�mQ
��{�=>�0c�E�� O^C��O��5�2��ӛ�m�ҹ�ޚ�J�j�E �;�h�G�4T��)�J�����S:y����_@J4'��- ��g�g($��a]'T����l�W8����Y>A���7U�U!���a�O���aS�Y��6�����Z�4��1�+R�#�K�������H������߿^�GW���3���hl-&�:���w�N���>7����o��h��?h����2m߷?*:Cip	�Qiu��@�7��OG�7�]w���Km�g�7Sh܃��Č|���'�;���8��p��|�c��Ϲ���K��{��O�����[��[N�	,�Z[}��v�a�(�?�EjY����Q�_G�d����v��Z��گ�*�Z`����V�>#k/��+S��R��z\,A�0�<Z4ۅ=(�k�N,��8��G�Ws�6(�0��5M��^�*e{	�w�C�ҾMfզ�@�˅B� �b�B��x�(�LD���*�Sګ�5u��A<���f.�	�0.ƍ�������}��s[r4��]Ga����h�2�b�bS����=D��=��>�#p�<'+m����X��?��E�E�JdQ'k��/�����*�h�PP���*��]�}D#M��ȢV�9�_��f�W��
�/AɜT��R��nj�V�8��y�!5Ō�е�(��B6���K�%�:�D�8��b1����Ֆ
����;���<f����v|�(�u�	�Ǥ_09!Mf\���������T�cZ� ��������t������Q������[h4#q> ,�)����l�71 n���n�X��6d�;���ʄ=+D�$2��؍)JZ���r���+��-8�LX1����EX�QI�18i�� f��l1����#��U�L53�0_h���R�,ʀ��sɾ��i�T%��&�b@;��Z��x�!9X��;�L�|n�J�@��h$O=�韏!V��p����wνdjME���>P�6n�um,f��L�!,���]~ܟ���ZJ����'}0)����Y���t�Lr	�'�OD�c��@�&d&�����M��-����4)������Z�JԿ�$���Hd���� �����f��h��w 'z�Q�ݓL0���&[_#�ز�ߤzw���Y�	�����m'��H�_ 0'��:���#��~��A90TW��}I�_�v������In��%ԭS;�aаy���ߌ��QqG=�Unی�;rZ�KH3Mhz<#z:4����t��d.7&�m[A��
w� m�{%C�&=`����f[�k�zs�Vdm��Of��b�PCʨ�����<�c�S�����}�	�j�(�	^����@D���b%��86w�Z���8��Zœ �~�P���Ĩk�"�M�ƦV2WK{���w(DU�\t�����AC���,
1��7�pK��>�������^�%/u�q�WH!~��$��@H9��ҁ�~7F��T�N��J!*������^�s��4+m���珝a2j\'�_��6�f���#ݿ|��.����=�̻�o�-<)+`���$�8Hu4�����7I���jV��������ޚoJl6�c�1�E~b�������f������5�!���Ug�ŉ
�N^�ѥ����	L������3I�FH��ۋ���Y�4@7�3�!��C�+��*�?)��/�dH��L�~�`��Ѵ~s}'b=�ɽ��L��G �F\ʚ\��'�v��e�����o����f��������S˙)z� ��o�mب��W[�s���c���f�\]��Τ���[$-�pF	�q�S�|~.B�&+P]��vWr#P7ƘSc�b��������X��#U�W$#��zG
{N�\"��[��!�P����ӽ�T�%8�8 ��	x W�����Z�8jg�D��΀L����'��-�VW��}y����e��/%/�!�|�7��+)�v�T��l��R<���^}b�A�J��
K{�p=�H��j(OJ��pޯ���j6��y��.��Z�c��e�Po�C�������H�@އ��l�u"�sS�Et1	��
��"�67ϡ�ԠKa.�9�ݣ�}��N��B�i�����L�`�߆!�$A�T�U��;����D���3����<������]��o��Lt>�{����/�<���<��╯qm=F�J�pv��iŎʷ�\�644ķ�wJ/�߬�����|�^��P9Go���^x�A[���Q�#����ch]�k�������}�w��*1=$�^P@1�YĴ���/��6�)SyX�n�	3%�t=�d�o
�d��Pk�LV�H1����[Ч3�F  z)QnC�jE�2��0aHO��nc���έZSrkh^�!��t@�ǝ2rDY�5ڋ�D�Dl9=���6�՟��U�h2��|�P]�f��$�w4V�HxP�P�Ut[�Ն.�w�
����?���0���Ty�枖���3�"�I�>�s�����IT��3�N�����Y_P�e�'��e�J%P��}4�[����MQc�����2�����2:I O�r�7��KK�����P�9���(��ߗ=�9�;bL��%7#��b��v3>F����a��X�:�1i}ض=6HA�b�;!�g��M�x�e��D
.����#Pl�;�d�Y����{ԡ�gp�P�����}�5����� 	Rq��I����p�*�0�������G�k|�M�mn����]��AVtO�]�p�"ēZؾ���3=�f2���~�~��L���r��&ۢ���=ٍ�
�Mt9M�Շ�$U�2_E���C����xZA���`3R���{U�%:�b~��}U���-;����6���b��� u�q�m,�����t�
;5R=)��[{��m�c �����҅���)j.�N��U�H��� 81�^X��o}}�!s̝��H�@�۪���31�J�w��n��SvH��zy�;!��:�i�Z>,�(>�R7��y�i�G5��z�sD�� Ԗ��4d��R�75�M!�E�k:��l�Ω����3��L|4߷���p�CL3��(�r��-7c�L,l�)�Џ^�j'��3�܀P��$+q�v: )>DO�ÿ�ٚ�C�i	Ͱ{XO��:,�t�P��;y�k�4���!�)Ay@��:cOO�R>�Ҫ�s������3 .*k�xf�clxgF���eF��W|��,Uٰ?B�g�eg���\t���H�MAQ ��j(ӏ�[s}Z��@�������?���9�r,�]?&<)j��#��ߥ�A�L���>�\J�JrT��9�Xk���	
��"$�>i(R��h��:VO��LS?Z�e����|�c�kG��1�D�t��Z=����jE���d���-�us�R�
(�,$�]XJR��4�K{�1��Y	f�;.���NϺ���
���M.���p�����W���xP ��x�T:����O��)I_�s =�R�%�aC��G�7�������o�L� ^k_7�`'�޷�'�2s ��ߢ6��ű?fUP��d��am-�Wxd��GU��m�/���G}O���<=�Of�m��v�g�S��<rֆ(�K�3���̋�ek���5�fD^7������1��Wx.���؟jK�+X����Pų�3�ej	�W��i���^��>�N�QW�>t�i�7r��!Dj��nG���J��^�g���m �>�f�� ;?�[�W�i�g"H؞�Pa�Ú"h$׆b�Y�K��ir}C��i��©Ň������JmqЋ>iH��of�\;����e}1L�������MQ\�ۏ���d^,w��c)��5��cg��e��Q�@�?��>~]���F�ՊDS�&)�0��(-��mS�و�����|�����.Z^��������gi8�u�8q��'`h�K6wo0�)][T�qn�����㶗'�Muw�V?��@�l���qg�l?�zY.^�~�8in*a]�x������N_�lj.��p~׃��JR]1�A{�/J�;�ޛ��}�KgFt�x�%�p���0[0� ;76�|���t�P���Xc�8��.�Ѓ��i��{ae���m���sؕ��d�R�AF˄ȭ�㋬��bc�a���A��}3������r�g��xx%~�˕c�ت6@�%וX�ᇭ4q�oL���j�C��x*5����΋�ݏM@F�/�ϽZ�9��Y;LGK�=aO	>��5�3hs��.�Ѝ����gMOx!]��=ِ�݈1N�P����}�a;��еq�����{�؍�ǂ�J�E1.@�|�{!r������o>�1�׎�e ��7�X��C��]�q%7LSs���lX�nL69%��گ����hźL�_�sn�1q���&�L�e��W�MV��{��Zqd�פ�w�֣�z�AHD�>_��d���������E�Hi�@�	bɾ���u�<Ǧ�H�~�����9��l��QG���m���%Ձ^��+^0�l_�`���AO� ��8����;P�Mu'��egƟ�Z�	鏦�S����[�:�A9Hw�b2?"h���K�k��-�	C�l�/e5%���K���
��OH�B8׷��<�͔*����_�:T/��ռ�s�:e�Yީ���_���╽�Z���+f�i�17nUP<����9�φ�f�/�z���Xqb��*G��t���ݍ��칒,�z��2�O$�%;\Y*��e��M���%�d���(�ζN��\&[N9Q���b�-ph�}�!~/��Mo��T�:U�FҸ�Jb*�Wsb��_O��a)�=�ڌ��l��.J&�Te@U"�e��� Dr����M��Y ���¢�w�à_~~o�y��=�w|S���ep^nb��'h�T��1�����x(L�-*)����(_ADV��A����0>�����d�zX���sp�i���aa����+g��o�Bv���}H!�R������
-c�� �R���[k앉�~H���&��*��+��G�Y(0�)���m���#��q�T�doЎ[�q�<{��+�G����(�[l� �)e*oxK#WOX�"�&_8(�ټ���zi�YH�V`���њ�0����c>�A�]�h����u'Q!�%��A��tk%J�X�{=�ҷt�E"���ښ�+X�� S{bՏ�3E�F�2ٜ�P+VR�����$΃���g����}�I��f���̗����LwZ�е*�#V�t�x��!w��m�ɺ��j��Q�J�����h1d�ZĒò����ب��ֈ��[�
���-��
��k�3B}!cOV���(��O?�V,VYBWm�a�W���c�KƄ��Gв�_��$�ey�N��dD�/,Y�*��qh�O�l?L(<�S6.��b\�A�/fr$�E���klj�^/~�(�-g��2����&uyu�_X��B���y�+���h��gQ<?�ڞ���?L�e��r[�`�3thX���Fo�{�_-��s(�FZ�W����z% ��1�+'��B�?T�5v`M\ALL�/k�M鎦�fJ�TRi���S��~��Xؔ�-���W\�_��.�����&k��e�������0Ǹ��ӓ~����ƥt�ׇwm��w�[�ba���k6J�YJA�Ǧ��A�U[��Ό8Z]�4z��	�b}I�~Q�r��FI`�����͖$��b�{��K�hҡ	��y`��C[�:��e���p�v�l@��0�:I��NL"l�i8e�� ����m [�z�F������"�Q�{��.�_�C�Pg>m�̊���=z��,@�O�6��g&I�6��k��^�m�.�
ʕ��d�3W�ߔ1Gf�e��ڡ|��?�$s��+���x���n�,��?�T
�$�SL����G�ɥ��:aC҇oE|C����F
M�mXg�x�����[�e-�:ܗ]��\�|5�=�In�0����2�O>�tOJ�yɯ��G�)1������?��^�KHI�P߷�y��裙�¬���.o�`�[��xߴ\��j�|�Y����]����aŚY�u�������\�+�܈�ſ��;� �+�4�V*]v]!&�{���(K�gË]ߌm�(1�e0fވ�ڢ]z=�X)佥AB�q
Ly]'�?�Y��X8�B|3X"�|?{�+�L���� '� �{b�?�%%�+�Ϊ��qK%�e�*qw�Y@2L0'-�١*<�$��梕��hw^-LT�G���qJ��H�^�-4������R�j��H�m	eSng�O��U���>�"��r��1��i�x(�|A�������_;)�Ν�!U���ܨͳ7*�]��-$+Xj&��1���3��I����h���P�S���P���{Q��R�X���icI�)�l�	NȚ��}�n���]N��b!�Ծz�������Uc��iu����P/&��>_�G	)��m��h���,��_�'����O���N4�٧�~\�����_��1oۈ���_f�RR*	��-�2��z��08f<G}�]��rV:-fd�
���%�*�3x����Я#�N�&E�^5g���6����Wc� ����6�6�U^�ʂ<��VI�~�Y�.�$����������y�X��҂e��wq�W=ey�N錟z���Q�������$*���.�y1j�?
�����0����ވ�����)���[e����Bg[\PsxS���U	�Cv&W�N���wcR��.�d.�g�;$=�vh&R����o3F��yU�_�Jɨ�	h;lj۷U�V�7R��f����4"�)c�v�Pj/_���*�œ�ԓb;H�_=�>�0;�[�Q�,*z��u��EU��lM��%u�%>P��h�x'���B�sb�*�s7������������^�E�צ[�o�����-"3���I��J�[�V�N�W�G���
HV��t��,`��^x��Q��/���bO��h�9C�"G�T�6�dRHo��or���Ģ�����~&I+���+�\�i$kvQ��C !w��_E���&Ҍ%��W!"��'Ƅ(Y�tiI�	�	�8����gә����Wrp�Kg��Ω�A��b�С�7�/�z�S9Vj�6�5+ӛ��=�1=��\AK�w�wx��ι5�~�h��U6�0L6g �)Y�J�wc��1Z�a���rn�,B֔�����ޢ���1([<��~C��σ2ɵi p\��E���4��rd^y�C���/���k�FY`	k�B���{h@�suL7�����	��g�"y�b����zP����=61�u���&�4��a6DGA|�έ�k����2�{8�M:��T��T����m����%K������SvE9�c��CQ/�t�G_�#��P����G�h��|��K�˼4d����~	v�����"[�'�Y/C'�s��e�&JI��M��)�Y��X�a�%�!��A ,�7~EE�_K��l��e�mR@C��m򷻝K.J�RN�bvG�G �D%S>�*^���ԝ��d�0����5�n3\.��h�	(	&�;��EMǋM���z^#����=ۅrN�Zc�A��2	��@I�s�+�z^��K1�����}l���;}�����]0|.m*�:'%I����ǰ�������Y�#�3t��Lu;��{W��vo�O�ul(u�g�6GS�O���˗��J��@�g�� �.�U	��?�R0D�薗� �g�f���i0b�l�G��'{�}t��|A-茲j!��b�>޺y��[|
���H2Џ<����^�_���V��Z;_���:�J���kz);���������{!	��O�^]���Ɩ���<+l(���;�b��!��������%^+��!�`JD�(�YT49�x�����~V��o?F���S.�Hg��I!��q6�:z�YH���ǽ����L ���ߚ��7�=������X�y�1��/hI�z.An�����j$���F��4�+G��=y}_�γ����,���#CT�br���I*���t��C=��[Ӕ�@��"0�@��sf���S���ޜ�P��=h�H:/��|Hj5�Ԏ �\��_͛��aE�@H��M�
����|�AF��Q�����t���}�p��~���ǁ�n~#�"�Wl���T���&6���ݭrJ�B0�øWŸ9�4h:uz+��)��4X:i:i�ni�0j�
��+��|�eLѧ�C�)V�'e��'t\^qh鞕`�7�נ�j�f(�����fm̭�X��eq����< ��0a�s�-�S1��N�
��9�܁���m�&������['��q	���3L�
�~7��R}�A0lȒM�!�=F%dˏ�!3�Q��/]�1͓s�|�	��.r�&m�:�4�w�
��i9�Ao5Y/��X�tu��䕙M\XKi�I267₇��7�*�W6�K�S�o�ɀ��p���P�ӵu�?���9���ú3摃,)]�Xc�)Ne:���Zo���9FP�c���ߒ��$/��5�gIDkh��{å��t��et�\�~4�~ǁ����2p�o)��T4��0IfZ?V¶: @���ݒ0�f>��#~}��my�J����2]�P=J��&�c~A.d���B)��T��J%N�("H��}��6B�ߤIД!��K?�A�È^.��~�������b���� +�e�c����H�^�3Zְ���2��3Hq�E�u�>a����1���8�~���õ�^�z��{�¡`�&���외��ObG�v�y@�4 �<ܫ��$�@���J��dgMuD�?ޅ;�$C,f�?kt��Z� �����-ۇo 5Fy"
CcG�Ю��O�&acrp4�x�4Ծ��I����D3ix%���@]	ke���X,v����n⠄��ˬ�]&��m?[�i�����A�Î)#إ� [�dZU���8_�-ޅ���n��jX��BhB,W;��=Łcg�7J���-L�2�$7�9o�z�$���S��0�w����	-À&��͊	q#Ų�ZՒ~F���
��2�FN�E5�rIe�w3k����1����b��r��<1!�G|�х&�Z��g%׆|	B�y�1���.ݲ��7r]�|����Y�Đȗ@�g��0lR��������l�R��)�T0�t��B��hڽW8T��%F���VH_Da�������{-�K>H8bX���0U�'Ǩ!$��7Ԉ��+�*R
�&�O���Yt*.U����5������?:�^X�Ӷy菨�jly7�z!�;v)󲔇k	�_	|�s��d�x�j0�'R�4��{[	��L�/��h��*9 �?" ��x(�ۏ�`��^;|��ј�u��b��w��t(P���_.���AI��
�ZԷL\��T~� ��+oLL�.�Z��V�%{����ܫ9
����\�����f7@��=U�cte��aE�<(����J����/d����h����Mњ�=�����(��J�~6�'�j X}:P�Պ�%J�M7���[P�=�'������]��q��Ί��T�v���;�c?�����B`߽�Dk�r��cZ ����� �ev��K���ʫ��6��`�Kw�9G��#�SY9��쫤R2P�����w/��a�?ܒ�,���LrKuN�U�������o�vKa��-T�O$�ЭV������~�Ǻl�h~z�eH�q]�%�=��dq�oGH¶HrnW�������8�)n��2,-h_O�V������=i,��!#���P�A�򋯀�R��5�9~���A)�+��C>l��
�J���CD�-�M_r����I��s����p�߳s_��lo�)�Kۼw�z՚��oR�3�7�F|d����[)�$�m3:�u��RS#��!�"�<7�*�����ؚ�(�oo5�0l(�X.@���q�U�+����!g��7;W���pp/�u`�"�3�y�R]�&H�K!lxy4�,j��g>"���\�qH��s��粻V �$�c��Q��!*�xV�܎��~8���%�Q�M��{�L68&�)�����P��H>l��z����+����eA�B涉^a
6��G̍O�u%o�}��@v.R3 ���vj��&��x�y�#R��eh�XQ>��7i\�ݶ=B�e�b��ƺf�m�S�^�"3�:r�H^=��su������n�b��ٻ���E�[�d��Q��|R�]�������@�O(/AV��5�f��L�V��?�?	m2�JV9 ���x@:}�wb������H:m��u�o�<a�Fs�k_��/X�/7����7���ҡ���!Ao�_J?�¸x���7'���f|!=�J NS�9l���9�o���^e�$k~�[�p�e��`2-m�,!�A��*�zǰ�k�E�Oi��b��k�Y���O�}��l@�.Q�x�T7�7��ʘ��O+{_7ﻬ'�?�zP|PSb�����o�a���M��%ZС���j���$��rѢ.:'8�� ,����#��-�
�qe�D�����H�}�T���R�����������p4M�&�ji1���sP6O,��Ћ7�y�f&���- �rmj�V������>�3K�n���u�z�L�wUq֒B6�@�ε�3�b�t�2�N������z�o6#]E>�o� $t(�6$�r�����a��M���G��LC}?
\*a��NlU��@���������޾^,���I�O�USGW��!�����7��<��&�����Z�у~���8�]��;,�z=�9��\Do���{����� [yvhwu&X� >��g��������9T�2�i��"���W��t��W��Z��w����I�/ti;s�TR�UnX���x&�Mڌ������u���/�4e�:��)Xl�6D�c8��#��LX��z/����<�62����N���Z�8)��I����NF'�U�k��,�?��
��`.��{�.�KB�{n��M��"D�n�K���L���T�l��NϺ-��u��)M�,�����_mK���A�K�0��Ԣ�W��S">�����)�x'u���5�I+(7��:1�b?�E�W��r���8?r=����ʊ�ߚ���~Z��KS����c��j�!K''O��y�s�[e�
Y���K�"yDAU�_� ��Vw����Ub\Y�$�͈�-���OH�y����>���|��iʭ9=W�c ����<LC��8m��C�����9��0L���.�<�,�_�LӇ������ەv��8�r�j�<�8j5�����3"��%c��\lCķ���(�zo:W�-�rr|���NV�'5T/P<`��Ja�$O������_�*�)x��r�<�3�$��\wy?�\��P62��n���aK��<R����R�5l%�a8&o�׾�G��M��''DBZ'��2�g�;�>\%��-J�5��.�\�A��K�s��N�x��ntR@'�<����حk�:j�|�-m?�Nps,Bx�x��I���T������*mg��~5��))"Ջ&�v��"e�$-.����Yf�aNb�G������={%"�Y/���)v�v���v.7	ӏ{��-R;���^��Z�H	����&YB�u>�
�~�d�]h��'��Y9R���>�*l�;@���s�U�F-��d�S��$ �5��Vv���U1�:<k����w��e*(����ِ����&#�Z��4e82J�+p*�v>	������d�p[S�'���:�SB2�\-�.���|�zq���{�(}�'#�y��m�=���6�:�#��m\�" tth���"j�%��U�蕏�`p��x�(�Ga����ɏ����-�"J	��ڀ<�t��{�H��������PX>PCf6p�d-�r��j%m�tm4=��u��J`	�#�����kj^����=#�wVT��5���c���6�p	n�'9�"B��<sV5�z�Fŵ�����ЛK��#�K�?�`G��£�n��� )�?�9�D$2?��YG\�$T���G�ؓ��}6�v~�a���b���*Z��NM�"y
��r�$3w��R:��p7ĢFF�$��Tx"!�����c4�����W�jragg�?���a��!/ ��L�s�� <���[=�߱��_G�Tf���rY;�'3��l�E�,��s�
bq)�Ź��aH��A��:�R�!O��y�& N�?Ʈ������e�� �H<��v�	#/��O� ��_f����9��2�1(�C�%Odz����2ޣ�����w�3����bBe#�`_�<8���xw �9+G��J�n=�y��6����<�Z����5&e�k�m���HNl��7��5��cP|��&�Z����8�pg_�g>J���U�ֲvڊ�+�~,-c�ßMy�%%W�dᧆ_je�fS� �̛��1���G�nۏߡ�Ǟ�#�����j�RJ�U�qn�+�]�?d�l�-X����i�z���׏뵆`,J��t<.K|�X�bU��� �8r�2�� �)9j)Om4C"pq����3�gˇ��?�4e巨��/s��u�SϥԆ&`��9�u��bt$-�vF}�'��Կ����o���.T�q�m�7x�	�H�� cҋ��4��z2!�XF��&�%��^ V'
���-.�'L� �6�ݟ9Ǣ����sY�I+N[_�"�n��ޤ�#��x6<����)�}�V V
��������q�|��%�h���ū�Õ ��u��W�� �C�.�0.��27�X����-lڰ����5��۰a*,9Tn�`la>_�JL��0zSkqM��q�ș�aY���5ҩ��.��ݘ�.^�^:��|G�������|C���!8�6��?J|�Y�����X�ϙR Z`��ʥEC�}�]�q?��`���I'-z_G��q�Yi��}����4u��b���\�@�� Pz��z��r{>cdM��I���uM���t��WAUr| M ��"9����w�H0����x!V5���{hF�ʱ�>hT��r1�Z<	3cT��A��z���#H�������;��V4����Kn]�(�[*2o����H��ǕOa���e���b�B�kg�M�5yw\b0��k@'��`/"�Y�DSo�5��n���_�9�*��m��#���&�83��i׶��h�&˟�2�S��-i���4ک�#��tk�&V��`B�GקN��ؗ�����| hD��8"�>I�wɩ8�J$<H������H��X��4!V�6]���%�W���Vt��B��!�.��(jȖ�J�~�b�	;�Vc ����f�B�g4ѹ��G�6u�s� �"A�Sbjy��,QE�k%]b6|�����10�����A��Ѱc�F���\��=n:I��N~�A���X���o��Q��̶���=�t����Wc��?�Աc�j��c��>����X���� /���U\S����	Oؖ�~L�ǆʱ��B�J|��@�T�FW��ma&�n4K�P��2�d7��=U�����fzN�V6ڧ�]w,7�|Ldt�/A1����C2�l�$�d�l����)��3Ef�1S�5���{�۝��#��Oι!�@�t�$B������Gk����'9ӛI6g��0$j�������	W9��eb�K+�\�Ԋ�m�^ϱ���q7�I{@?�"��1���$7S���ו��c����кid�ARݦ��I���X~�1�/�{O�+'r­T���c8ZF���mO^�_Yj=��"Q	��C-���o<�St�	>l���W&�8hV�]GCp=� 7�^��]�(�^�{y�#����)s�-��<�Uҽr��V���"��.��F���0�LL������r���W��*��D~A����\������"f��]`�(��Gh��_Bu�M�n�
`gdl��#�?2��S���'�dW]>�X��7]H=�l頞�˞�?� mP�s4u��;���J!68�!������S���61�
YVXY�,]ƹތ�:��!hY����?~	���>S�3A�62V���MYC��Ske��������݇�=�Y��ϋQ:3�~��"ӢU�̜$�m��Ж!u�CJ/ �͚�]�L1�kX'������<a�p�O3�>t�p0�����5+���V1�����r��8��&��� 0�y��x|}��b�k��6�b�6�o��kz
,��X�Z��������J���ɸ٭ph-�d��v�Q�s��漓���/
y5���y�7�&a�_���6�8
��p��-��w��H�e�X��� ��y���!�X�C�R*�W��:����&d�����</�?�vνQ���:7�������F����2�#�������0_�����<�[s��["�K-�����s�k�'�������gŢ!Ȭ}�q�,�XE��2]�QF��''K�ܩ�����B;)�܉'^O��Y�������6�4�e<�OGG_���/����?=D��ҝ#=����8F	�Np�(H���<����#�"�&����u�����T�����g�u.0Z#	 �<�t�SX�Y|2�}���I�48YS��+i�Fh��E�Bλ%�U�i���)���7Gz��cqf ����c�x+��J�C�J��0h5��POz���vG�ۯ�?ɨt����W���F~)Sʍ�/�_sȹ,X~Պ�e/�=PùP�]�d�U�/�O})޳���3�^bj�\q�w�ʆ|�-_Po����*U�P[�uR��ʑ(�\��[9sF��PR��o�i�k>�f��I�	����3h���-�j?NN��`�J��j.G��עŝ������:y���Ǜ��峈��[�]��j!�s�y�§C=k���[���1a�\���,�t���j��EN�����:;ޜf�Tv� c/��n�Ǵ%z砝�_k�������-} +E�l��֙-�aI D���$�r��k��ˣ�F�6W��m�E4/�3�ҵ7C�0J,��"y }�Ҋ��Z2$ds�s�rV;��i+ŕ�5��^$� �Y�I���0So��v�\���<Uk�(JJ'�>��χ�����V������&��?�bq*�h*���L�O�xP*N�[�n�bsy���x��/�4L�]J{{*,���5�O狥k�~@��{Rk�y�f���};E;��;(��j{���]���<��L	��Wt���
�}؂�,޾_#�s������h#�#I	
��R��@�?.�"�9l@�X��G9h��|�}��y�I���)/�� }5ԚW�i4�E>���ns蔲�{Nmr��~��_;�`���Y���T���*����?0��R��p�N/�U�|�K��Λ�m��J�C~�2~�X(E�����B�p�j����'Mi(�v�Jd�|�#^�fuP!g;ԍ�[�/$�i�qt�9E6��&Vj��EtHrB8����tR�vaZ�������V�p�rL�ki��磕(x{۵x>����IX#ư�V��w��{z7��4�ue�|:I�����ʛ �ed[�r�uaѮ*�p�ax�=0�R�N�;�8.��X_�_3Oz���I4�aV�����@޲����B��q,7C볥����c���$l��,���~�-�d�P�G}x��&�ߩ�?r���E߀�'�g��~1C�����2Y�+Ê��F�A��ޓ�Y�Y�ЦwF�Z.���Jq�?<�Ee��(LA7�ɟ��M���R�;T������� ����C	�+�=�Qg�J����w:;��1�������-sq�5����*���@��w�w�u���E�}j�q��W���vn������]��������*sT�&7���m��
�J�?�����V'��+��/�mFcԴ>]�{Q����h.�q��ci�L�="�߫fT��f��X�cT�>�y�V���%8���ڜv]G��eA:5�����BF�a�'ip��)HYUT��w��]���E�]k�H�'h��d���;��0��/�f:Q�� �_Ly���c��Nz�tT�7�bߍ9����o�ä8n7ۭ|ʚ�5�}e�&�Y��bZ���/� _�1�����	b5w2}�EV�~ݤ�����/�z����Z��
Eq��x)U�xt��-טVy�/�#p�J;!Y��'�d�3XWgq�|/r~4�k� �N�-����밓�lS��y�H���<!��.VI��=NE鶒��\nA���|�1@�± ;���(�/ª���6BT�WGO��N(�.sl����z��>����b(|�i��#݋����:�f��r������ႁtaf-�4��T�ځ%�9ˑ0',\V.��5����<�~Nb�Ro�Sπ}e�Ė/�~�<$����i�QԶ�k�#̶��e����}�&��e�(��P݋�q�|�Q���9W����A��6��S�]y2��_���^f{i?b��2B���X�� �'(
�e���+�G�	ȓl��x`�^bO;{��	��O����z����;vGe�շ��s$5�z�d�H�������s��X5V�Y�s���>�,h�q5�{Aۭ���h�$-r��c��\|�|�у��z�����vt|�
0��j?+��QA��"��Ƽ=����n���E'�SJ��/��v
�#��u��%3?/#!ز�Zէ�k���;v�1��:��B\Wa�S�"���_l�>��<�1A~�ڑ��Sfc���Y��ˊqd�,�o�3;�I԰{�4TRF����\��M0.(�긥.�=��G~v8w�:�ᯏ[�k&k�m��kA��{_��(����(;)>].)Q,*��T3�A�`Dŗ`,�T���i:��+R{��ƴ�`���M�'��/��Og��a@K���B,�$�C%�ܹ�+����@�I��Q�n_?�,��!�Ov$]]�`�"�	S�\v�͎�eN��<njѷ��|R��l+Mߌᛆ�t�V�H8��U�Ja�Sk^/���a�	ܹ�3h��A� ���j$�1*&8�	�O��P�E��/�8��HR�
��I��dT	�u&�I��T��Ї��vU/t�1���2;v�����6
�w�s����&D9�7���Sƌ5'w)�_q�#�gr������Y�������L��R��`t{l�_~V��SuWϐ�L�.��۲�l�L�+ˆ!p��i4���=��+r!}R��'>/� ��ۤ���	ۓ�Z������ki����%R�0Τ�x�o����\��g�'%�����p�5T6(�0eQ
��ҝZO���K��z��yn&'�B.�s��#���j�=f�� �ݦS��y�
��0����M'{]�@��z���=::_;S���ds烖T��Ge�Q7�o����5Z�~�Re�OnQ|9�cd�3\w$�.!�	����ƣ����t����ݛ3�\��|:e�Ƴ��UVKHؠ'��t�(��]B9:�YuY�%�=�|�
ޜ�7���AYv~��eң-�z���R�c���z�[�%��~J�6a�k�{hf6�A{�i��=	�:{y�����'oԬfe�P)���q�^g0�#Qm��B)=�¹NW�$:�2�� o�O��4L��6{	)^��.��Lߺ{ܵY��������6T�����I��]�u�l� s�|��V�	0�:p� ԉ���X��4�
�?�Y
�3|�M=_ϒ���7�gI��g0xk��_���ӥ�i�����T��KFA�8�4�9�Ľ 	�F��v�1.�F�h:�&�6�R`ɷ���Ph�|}V]�y�C��'+�rR�{�ވ���]u	�=�f������:VUz���Vwwj)�",n���dp#����k�N�Gp)T� J�j�0���KcA���;��Ӕ7/S�]x�k%\ÿ<`~k�� �������S�4k��83��OZ���U�[۪��� �K2u'�����:6�=�.�J��5�GV$	�����^�
�e7�}��ju�[�S�}�����S�m�!FsdvY ��b<��!uh�]f��O���8Ҳ���G��9Euf����VZ�y7aOIn){- �xC�Z<9�5V��)5��fӆ��q9��LL�P^B���i[��Mv+�nܝ����}���ɵ��UY(g��G��K�b+(ی���Pd	0��ۑ�'���h�� ��^�Lxq�� �N������m@�f��Bw���B]�߶E��g�7�m_���w^�ꤿ��:�e�U�����(�'?p��x��s$����~�o��m�m�k�#M��Z��2*�?�#�h�}��j��`Y�SU�v�i[����|ڬph�V��ÅMƎq]7��+?�Ӝ�${u��1�#�\�ᤖN�w/Ծ@�ic� ��vL6���$�R��t��;mЖ������H�rL:#��XMf��7k<���\~��qP%�	g࿔��L=V��L��v�#5�+`�d�\�X�$�2�����ɇ34���g�	.��T���d>��w:���#n�Y�R��K|��-��ɜ5�+����\��UY~���4|an�_3�r��u�(v+O�3g�e~���ל��c���n�c�j��^g�]�F�^��Q�k���<�YHȇ����)4)Q��LK��C�;�>"$��{BGF++��$x����]L$~�f�{�&n
֐z}a�d���N���*�AO"�)�� E��H�K��V�N��=��
m@���Y�nv걚�.�N�S)�p�!.a2]�B�8y�2b�j��*%n��/����nGj���EH,��_���hY��y�A�Z�TZ����c�����|��N
��ش��xEJ���.���A�4*4��,BQ2줮S� �8Uv�O�yxm^7S�@�����/��0����Q���O�	?ҏWi�";LHj�
'�*+Ǧ=5{���O�Mǚ�2��Y�ش��X5Vk��Z��.�Ϗfv����B�x��φT資Q� ܋L�K���xf�%��&ᝫV;sn����*v��rs�×����`5)B(Y<M�2aSoW��M�z7�S�m�
M��m��FT`-Zѭ���=�R�ò�����I�8�
�dT�8�s�7`԰ ����J:�Zux�r�¹2m��
�܅��(�ަ��������33��U4?�\
}��HM=��YONCڸe�^'=�'�0�P���94p�A�=�}USĊ��b?W2��C��ڦ�?*�OE�C�u�@[�U1�u�ҵ*(US>���7S�!r��˕�u��?���닲��f��S�ijs�៭d=1ǯ���%�٭�?^��*C�tbJ[s�e��Wï�Qss-��A�����u@�����t7�Y���LJ�bS��".���)��#=j�����nm�W��0�s��1ǳ`���+��r����M�o�4C#'C:�MC�c��^��F�����`�h�o}V@�I�y�m�mzK0<% CSnm3	%\����L��-�(o<��������݅�3q��#Տ>k�f\/CA���/��r&X�����ܮߋ�Ǆ�QC��	�|n^鏨��Je�h�xY=��_�v�)�i��	o�A�I�1�B/�K��ۻ��n@��ۀ���BTV�l 2Z>�v�H�n<uǜ���nHa=��r'}�����>n�3GT�$?皌7�� 9sU��P��BKlbcX��.������6{(��d[|1�ݮ�V���W�0~��wK�̴`�uAA ��W�	Z�࿷��^���wȽִO�۪�,}�5y�P���Lփ���+&6RBخ��v[G�[�T�\5u&�͖Sԑ�;G�Qk�&���T��*�G#әs�Ս�.�x�neKQ2�u�bc�F	w����%_7�[�l-�!�S�lL4Q:-w|N��`#Y�b6����x�ɇ�n⃛�2F�5��ކ=��b�yp~U��9��1M�k�T��� �1d����v���>�b�<�}���ᓺ:H�P_���mB�kB�ĉ�
�z�V)?�W$'�/8C=��`�K�J�����{�**&r�����`�*jQF�i�o��Z��;M�-����>��R�V"�������髈�d]�p���N�ŵ�%=��3�K���1���M��|��#ߓ(�:�%S�n1�nj> )���d��Ś������h�(�r��s�ZJ�_��0U�pj�v���D3񐒥���3+����N�2���`���-�q�����{M��\���5�l�Ʀ	�Qs3)�_�ls�̺��/a�t�,e{6��ד�P��L<`}�C8
�l}��2=G:O�%�_��a�~�4�ǃa�������KE��[�o�X�j�a�� ��:���plNt�^i2��ޟ���w��"Z=�Ht!Z&6Ս�l�˞?��j��U����sT�g҂>��3ַ_��($[�S�
��	�x7�+�� �K�U`�F��\=]�rY���j��t"P���7!͈J�63���j��>�?���$c�!a��ժ�	��4���������0+2�rM
tw���x��]�4T��V�L�P�
���\��|u���E4���&f��E�&[��ƛ��7�VĆoFk��Cc�:y.���������Q���	",X�fJ�=��{r�����e����E����>������%Y�Zd�3X��xРϫ�?'qF,^E��/��k\��婴3pFȼ30�f�.<%M�w�,U�[)b�K̏���86%d�j��8���������7'��z\K��?�fL>H�#&�9�(�'X��`Iq������.d���0���z7Μ�A�im&bL�T7K~#�F����^h�S���R$d-f�^���<�(79K�$�~L󒁜��� u������s��P��$����e��s�U �@,�ˇU��_կ�o��z�)���<�ap1θbȘN
��y&�5?�>=}cQFk@6���|t�i;n��C��~��1�ˣ����c2�cU��f�^R:~�!7���r�e�Y�8�-����+0tZ归����q苶i��S!
F�<��z�u�tk'��gI�eP���R�I�qk`4S�<���C�U_�L�Y#Cb�Jz1��e��3*�d�1/0�D�4���ug���J�C �\�d�?f�Ӓ0�,��D����l�+DM<.�X�l80Q�X#�|�.�w0�C�?r�4�58��B
Ἷ�p�+P�w򫶁�� �c9��m��7bT��;rnLF�~�����ҥ�vh���-�ϑ�&�l1�1�H�N6�N�@�,��m;x���d�KLգ�][Α(��Sd���F�E�Z��s8m�ޏ;d��<ī:T`��4�0.!>�
�߸{���G���&��]�]��V��c��B/�ב{���M�q1�=X�3���I�k�.)M9׮�DC�5�c���>a��5���-[�,���A�˂�1H��:ͤ�(�-����Θ��%�h+n0yb.��:X7 z�A$*sK�~G���O���J�w�Dt:$�����ÓsG3bO[0&���h�D_�@��Ӥm�F��K?��W���)����-��Q�-M9�Va��!%_'	o�{�H�� RL.�62*�"d\nA)-I���}��^K�Jb@w�`�J��9�ֆ�����h�fL�k���&��d���/8�v:,�Ij����33����js����b�e|��ʩ򆘕!c���I�x6 +�~���o�����x����H��Ckr}��f��K���hue���B�X��>�~��)�	z�ɔǸL�W��GX2X��M���1�&��u�^���7/�����]<�H c)�oR��I�6��S׊Fz���J䉄ȇ&��[�w�t�tfں>�:�����Z�#�@w�ʣ^%�����N2�>����q�W�ǰ�7eq*V4pI�c�oU]d�(*��^���/녊0��g��x[iD�R�i�.�8�"�<�������ܪ4ߒ��O�"�"<�qZ����s ��o���Jc�L7uf��R��������"�IV�S��tO)̫�����O��/tO7?/L�w�D: ֖�vt�G�x�S�L˓���;�"kϙ�����]����w�� �h����UAY�lk"���wHl�D������	k�y���O��U�z/�y4�9[ˠav3%w�~,G��=�"�卄�h<�F�bpS0S��<�+�O�����[���e�a���U켦y&�P�+@zn�6��yw���+Fי����4(���R�e�*��p���d}?$�����=����8�.�'��Vnqk-僚}̵aLUx^���;�.��$q#o�4d�t���Z@O�d0�ZjL2�&]��E\��t[C�I�3e+�?������!GA&���R�sgy�V	-2.r � �mu������� t_��Q�¬m 5�Pҍ���ׁ)�{�ENl��q1���Fd��j�� E�;x��Ic�B�1�ǖ dkraBe�ei�1��Y�o��
�$^�/z��}T���	�E�S֤��X'��B����e(;�uRU��A7��F��e�QM~�Yz�;�o��f|�2����.�c���6j+X�t������*��[>ޘEA���ɕ�_�p������Q�SUG���L�߼a-�m�Ł �m���;�G��+���B5I*�ty[큐�����<>몏Pw�ݷ|�lo4C���Nc�xRM�B<$��qg�pYa�����%|�T�S��zj±�1p}��ΐ�<��������F9<���ǲ�)�B��bX,����8�+��AT#^��֞��Y�h�֔�9<���2�ٺ=�o|Y��ʒ^�V��{��v�tw�ڑJ5T)����k4�Dq1�۩ �F�l �7뤌Rf���*Gd���v���)�烘��=ʚ����ҥPQV�����)�=��}��)w���̝'K��}�]]�ɸ�նsoi�4�O*�-k��o�<'���zd��5m����{O޲+Su	���s�?=$ ���b���fH0�Hm��#�>:-t_�ρb�FvHRF�#@g�,��h�'���"�<�r#1#����,0��/xF�s[�A:���P/����$륤|߽��<���RoWgi�4�~�
�*Q����R��7�݀OH�	s�!Tˠ�
ӱ�KL��Ś�����%�oKFݕ؄�D�>��7��|���C�+i=���:]�ZH[��ȳ���^���e��I���t317�o^���AiX���N�� �x����u,K�[8���y�@����7M��=�⷏8�|�=��c4%��}0e����Z�kT)��v���1�!�+��#���J���HuT(P�Ќ�SJv���_��Y�V����=�=]�cƿW���5 ��-x�:1@��Bݞ��|"�OL0\s�VIb�j������]�A��=�ȠQ�H)��\x�H5 �$����7���5X�;�B�,{�$Gpz~Z] ����rzƠ�㷍����)�p�6��RuGXR��~��[pkgȎ�S�;Z�g�����������`]9���jX"��j&J�*i���i��3މJŔ��,z�� 0�#���Q6q�B~f�څ,')�A@�X��d���E����,��9�j���ZH�5rw���=bs��J</���v�=;���v�e�Ӝw�C�,r��$��x��9/�-��+Q�U�+�jկ}��d�v##��7�/�k)�c5��ΰ#sgv�� ������=,N�~���[	@3��$�M�!��|��$BT)�ئ*2�5�9�g�5rx#8��WE6��Yf��uWLSc�� ��c穾9qU�,v�ڔ�!�Z�ގ�S.y-���q}޽cy���PA�rޅp�u�r��{PT�˓�ܖm�9�����%����ܝ�*3+9��ߜ]	Xe̼��|�p44��а%��*
C!l�&4�VQ:���u!��F�m�/C(!e���K������^@� YKt2a�Vw��*S����%�;]8���<Pv{�7��Z�n����Fa�[�"���J���f�:�x�n{D�dVb�~.xL9��*�E�����Կ^$.�k��O2֊�i�eZ�����V����Nk/Iv���c4Ջ��4�J��B����������
�s�LDlSf���O��Y�w��	������iUG
�b�ɗ�6�#S3���I��D ��,�T�S��f��g3�_u�Ł�
��G�u��h�/K]�`ڕt�wg@�2��o>l�KZ�i�-oH��޷Z��&\�T�;�<oFX����9��b��S0��jB��xj��$8}˚�Z+I�q��d��ٛQwp�0��'tÈ�]�M���9�uw�L9�6�h9�A���9u볠Nf��m����wv�)h*�a���v��
�S�b���L�z�'պ~Y���m'ϲ�.���Qd�A@8�H͈��ٰ������Y&�恻/���L����ŅZ!�+tƹZ"v}gl}w���ۋES�V��]3�:r�hڸ�=�����T�%;p��;0 �.�g_6`eEX��|O��3�Q�kkA�`���x�+�L_�tA%�.��j�O�w�2��\v����x"�u�}/HJ:�Ng������D�:�8ѶY���a��Ɣ�n*��͑�0��+����'��Wf���!Q��~"�72�et������t"�of�؀n+� pW��/C��U(��F��pH'��h���{� 3mFg1���㿾m�+A/L�?jܣ���Њ������(�z��s���%uf�rŊ?��P��fA���29T%V�-� Vݦt��.yv��$a+�n�� ���`���=���SQ,NeA� Cgj��
�Ebn	P쫖���?A��������K=��F�<С�.K9��8��?��;A�z:b�Ł:]�)�+a+�P@Cy�Wy��ۉ��T4.��_26Lr�Y.p<rς�> ��X����aÎ;�����W3=�]@�oC�J��<E�fY�1z��YG�>%���֠�>\{�mt�bp���[=���.d�v^/� e�8<��CKbB�����P"H�� �l��7�����v�֮%����RvL��v�t8<$5ڷ��p��$���w�s��f��>��N:�\sL���&u��=�B�=�Q$��	�6Hā�	����)� d��>�]u��Y����qW�I��l�	4��<Y 6����B�9�O��9��7��]�.!�M.�Ui8+���q�	Ł����] `��ʻW��ת3D;���gq����eNZt4�z�:�y��u�h���,�S�t����z�=��o��!y�~PM�;:K,5�B�E�%P1�������K�"-N��2bZ�R�f��b�k��i��|�%o��z���P�Q��m�������+�����:6�r��e���H D�!z`!O��a�{v�Q/6�UqնթV�ڱ���+r)OH�?]Q��-{{K�A{�A�+��]7�C���{��2���{�H� ��E��mٓ`��U��b��H�m���~LT
��A�5K7ތ[�N#�	�6�������y�I��L�!��ҏ��vu0�TJ��we��l���w@�"q��<B��fT��\�#�R���?x>d����u�k5�����ZEIӵ������R��d�k_0���q�k�F4i��p�d�n�>�MR��N�OA��EV��Vd�Ԋ�7�p�ŀ�0����E����ܢ1��FE��r�a����Z���)J9��IµA�Cm�%1�����k����O��ѕ�`1h���-�͊�O�Ľ�6�=�������<�Q��T�6I����l�/aįo�V��%!X}����
��
>�ϑ��ڹT��u΄9z
��!$�C�����ӫC3M)�2	����s��YTO���EAV�u�� ��~"��qv�6�@͟���o���3���)xU��dI�f�N4/8J(�����ć�&U!!��Q���=�ef��`~,ZPÅY����
�R������vbןJy��2f��wH�C	G>XD�J��H������p#N_?&r��A���X;���g�T�ߤBI���|�9D����@>�%D��m��D_�ı�a P�Ѯ�k�i��x��&O~7�<Y��Ll��<J$6�d�"	��{\�&Z�D��Ar����Hy��FоB�)�� ~�)m�VY6���=��.ޯUK��@�Y��<�e	3jC�Y�琜
r�|4.�~׼��L�jx�����f�q��Uv�EG0
�1�mMЙX��ǰԞ��2���h�&����y2�<�ƾa�i�g����!$4@�yѢ:	�6���!��]�F�j<�n]C�߫z���ȃ�d$��](��*(���2#�F*{||�ec@lݠ�j�aǛQ�Z>��b��V�͙��J���*(f��D��ǒ�x���ڥY�2F�(B�����[���4e\h�]����9R���������:�����.i���,KPo���ҔQ�"��L�P�y6�9�u""�]�S������-|v�U�@��鍊��uo˹c��$t��?��e ���_-�K�x��B���Ë�H
�jr}|����8t�0{��4~��̳]
�o���Z���,�y��y��}��gJ~~.���n1�藷�4�\*�2NUF���/E5�P�"B�p�ʟ|�Dof�#e�Q:�G7U	�؆�VE�(��B�OIŬlI�d�t&Ka\.y�����l!챬�mf&�����VC]���x04�4ZF��z��C�|�]�Rŧ��
���k��˒e�:�?o�f/5w�����~m����	���C�+ζ����V5,�m�j��\�iVH`66Z{���]����}�5u-/������\0�|��V���m�|r��n~-8k/{q�� ��y"C���W��A��ې��{��:�
���^��l[�x#�Dܲ��w�)��춖l+��%	=.�N�bu��`%m3@yNo��P�]C*Ճh��]�m�J�B��<|ͬ��2A4x����
��5+$�<9�QaF�p06�nF�φ ��:�-[�kT�����ˣ8��Z+�Z��p�X@f�a3C�<�#%�{.cӜ�OG�K�"���Z(Mw���/��^y�!�/n'bm���j��F@�^����X]���x��w0`�u�±�r�}hQ�u���*�K��7��N��c2��b��B.6bU�[����!ƽ���D���5�]c4��~���zD�x��?�,�u$��~�.E��U;���L/	(�;z�9qrvxLh/�o���C{��u�Q�45],3ĸ��̈́��c�7�a.�$�4�l����&ߴ�]���.-��D�R�$W��"떃�GU������ز�H�B31Hc�Z�}��I�1Ip��#E����� C�e�o�?q�X9Sj��k&�Sq��$�g�u ��� 2fu�����fU���l/ �aF|�_�?Q����Wb�ب��+���-{ښ4�o7��(��e��<uTk��;���A�2��s?����k�f�#�wԕC�i�^,K��D�<���S��9����ɏ��_��;����k�b�Q�"_F-����k]���9�d_7����O4 �Ic'�~v��
Q����s|Ι���|���h� n���"��U��-�^��qI��B��ψ���9�RG�H�&�{	�W^��	U����OH-�o��"�{��J��q�����ǆ�j���,1 |��s1_e��G΅�-�d^����&������pjҎ���&V��\e��h~�9��N�9�O�,F�i(�J8��?k�qic�E�ѹ�"j����������<�HA���$ҔoHe��~�������E������N|OTV?a'X=X�Ga���閲�����e���]�|�^���r0?"���7�U$��<"�S�4m�L�5��VuLѹ���$��Z$����:d��� c���oeD��m��l�:��ȇ2��pB��c�2���1��%+����|��}�s\���9�$$-������������)	>�U�r��	e���^/����xE0���EϳMtU�0�'��,ih�� �h~`���N��x�o��~��m���ơ%��^m�C�t��y��a�HH�TȊ��YR�* �BH��f�ζ�B��ȷꬺ�<���?u�dN*/� /S�9���N�ԝ��46�>Ƀ`���.2�+��F��_<>I�J���a`[�����Zi�.*�vAJݒƆ��i ���!�rNHX'|����뙢KI�'�1�z��t��b��#D$�R6�ɀ�A)�pyOh/i+ج0�V%��{�<�?���qXL���a�iI �tsuτ{h�Ch>[S�m�|���
%U&e�BDw@߇�AH����:��x_ܝ�X�V��w���(A��K��N���Ы�&=.�}�7x��ܮ�(�U���~�M�O��|�ݝ�u�����	�h��
?��5ˏ��X�K�A���e�l�n�ͽb ���m2V��;Mb��N���,T��s�<�� �	<Go���)7�@�'�E�F:)o,=�Q�	[���|���$���� |q��s�������̈́�KU���\����{�u�M�F��G�@�fN�HA0�%���E�[J�(]�Wt�L��o?�����o���za�xb*�$"d�H*{�ʞ���d��Bj�w�sJ�13�x�p>C5�%�pa�Ԕ-*>��#�Ы�㤪�&8�UIt.��)���G���(D���Xh)X��X���T�V�=�ϣ�uWGo�f'U<z����/�qH�nQx;p'6ɬ�`�i�[�evd�4��������Gܡ�L1)T�YS��:;n�f�9~E�*=Hso�9�]K,WY��zL�����ڥ<�C���	xȅ�Y����͹\�R�R������ 1��s���UA�=+��(����>�::Og	"��g'm4.H�P���.�n|=��ْZ��B�>�uS3�xh��`��T?�~`�R�|U��4Dk��Al����'n�p8y�2��O}�/��&ˡ(m�s��zˉ�����C�Ju�˕i�62S	fH�x��]l�חK�ȹ~2B��F}�Gɣ���kkr�x��Ė�����8�'.1�o�Iݡ�ѭY6O&��\��l��b4�j=���R�H�A����D� M���\C�;�Z	��;�y��iü� �.E��r6b��S;���*��cq7�W�,2�QK1	"X?�����KC�c-�'�O�x�)��x�� �����2�D9�/�,��`r����c��]:x�>�G�5�]��(�t�rL�w;�F;/
'��j����n$eH�6q���-�x'먞o�ҏ#Dp�:�^B��(,ŝ���.y�U�d�_����O]���E|�Zc~,z2�)��5�Ӭ������ց��u>~8:�F4Z}�;�����l��{��(^uGt����F��~��2w�O�n1]{�Na�c�+�c���,�`/m���\� ;�g����U�PB�|����%Q2h^%2���t5f+rvێ���^xHa?A[q��R�����9�^p����`p��;��A��S9���]2Z���υ�4��pG���l2]<���o�q�7�B{���h�7�liƹcg�p6�������c8t�<�p}o:��uͿw<���n�#�޿؁ǣ��Ҍ�j>���`wf�*ZRNm�iN���� �2E5�
���O9�'�=I6
h�6���T��Wi����+	�'�q�o��r���t��h2�2f��n�mG�_�%�r�C�y��?d�;��Q�-I���%�E��r}*�	'A.Z��h�6[�1����E�,b5b���xb���V�2��ԥS9�Z����$ӯ9�V�֕x�I�l�0̻:w'����ɳ}�lo)�w��L���|�k�A�� f������$����Ю%z��CV���|�Lb���JJ1��2�5\�"�"Vj��z��NE>�$5�y�cJ�L7���9�ێ(/��]JdT��8R=Eëx�$��cz�e�Dp��ݯ��k,���:�� ��A_��I�V/��nI C^]Jr�9鐉��]w�q�iv���P�6h�K\�֓�&�їH���%e���s�q3	p��T�N�)��Ǳs�ۯφn<x�$�����L�'5�q9q]&�Ždk���������br��'9��G��U�ޚ6�2a���?�������t���?�\@�~���[��!��5��	F1о>�)�Zhԇ"w��	Lb�=?Ƕx��WԊ�v\R&$4E��?ؑxC^�Y;���k��QKֿ��I�� �]��>��K+�i ����^����0��ջ1s4�t�>MA��k'�8�wX&Ʌ�� Y�1l�&sZ�(��-��T0kĐ��3^W���:�U�P��6Ƈ�.�ɶ�`y�����<��{̈f�xm�}:��\�N���}��k1~�h��\����cp�Y��ۄ*��7�Ղ�X<��~a�5ˎꕥ�p�cE.��.)�V��
"�t��jV3@��{�Oc����i���+��^B���ܹf�&{���tޮ��/7�W�DR�cl){���y���2�����܊�r�7��Y�"e�e�|����W9R�Z͝T@+���N�2km����"Bs%��.	Z'��CI�#Y�,Y��IE�s���0�Jsǘ���b����e8����/�Ra�������43��~���I9�=Qp�)(�!����!�s�FW�?)IWkZ��9����ճ������jS'.и�L�_=�����U턖�6Q1֔o9=L�#z=�d:����s�L�y/������-S��v�ifT('���+7��dE:B^Y���/�qvó<��)��2��:�P��H�Y�}�7�ߛL��5jo�J�sP���1w灹ۛ@�2�X1��5.s������֭]��lq(���Xn�gɴ�RW���k���{GMey{|�fq")&���D�X�,���h+�U����U-|�o"IX<�c�E(��N�����@����1<�Q6���.>��g�{�%.5�Ε:�f�GdӔ��G&�9A�&ʈ�[�x��rL��\4_2Z+���=W�~`��s��,5(�e�v@��+�xq�i����1˔|7�W&�9'U�r�(��t��#5A�����i�E>%��;���;�� ��or�8Z3��슦a.?)�DR ��$6W�FH�U��W�"N�1⺮��A�gg���}�D�����A�t#B�C޿a�s�w,Tc��|�	��-M-��k�x�!��v�6gmiZ�1��mY��+h"�%��.��g��>�d*�:�:ő��%�����r����嵿���h"�%vgsH?;�P��
dG�=���bQ;UPר�6��s�V�z�#>+~��Y_]ks�CtU�,��6+sm��
�J'�_�8����7	��Yd������	E�w�<�4�#�3W-s�;{1&"��I�G�(ͭ�o}������S�i>�|[ϥhM��C�GgxD��2��=��_���,��2� f��
��ً���zb�ϸ�W�c��G$g���^���z�`a��2���I:g��N\��4������fot@i�c-���Y{{�I�r㡻�x��!��)�R���_�&�)�K�.O)��[��T�
CQL�q\;6�x�~�7d����&I��6���"�|p��׷G3�B����0&A�ayA��5E��(*���2֎"j��VЉ���m_�]^^��f�KR�Y|.�����b�S
��t��_�2H�҉m�g��D}�.G}"�ō�	�`L��&УQ����+э��~Z���hg�%��Wޞn;I�{��H#չ.�I��k��&��hW�]�!����uH��a!<j�exv@7!��4��i5������y������?�uw+)%�{?W����i�0&���t�H�	���z*/	��I�
����R�5U!b���j��`�d��W[?Z�5pdB�}'$�5���C�ͽ���ϧ��t���#k��S`TŨ:5m���a�Wl�
<L<\�ɘ���~:L�`��M������k���ƈ�<,B���^���x�%A]:�?�����S��6_M�J~|�s|�Cr��M4h�F��OB��!2����X�^$�ߜ�+#*ʲ���NBN�{՝*����msO4nZ�C����[��k6w��l�J����<|Qgh�����WF�kxp��ʰ����wS�c\����3�kC�I�H����Nϝ�ؙ��KF�H�A���?�+��ZE{��{�1Hj���>{���,h�R!@���G���u�&����0r�tZ��U�6U3v�F��ś�����I�C�{�7\��5
��G����Dȅ�o�8�4j���'Ep�|���D�z�ps����xl˹�)�97�@b
�'��;a�9Mc��4���;
��Y�ߧ ��}AEf[)ߕ�eo�,��7�1`�K����A�u7�Et���u/(�Eϒ���޻|�(Ea?Op�q��i/�H�ݽ��8�6���F��p-�i�
4E04տ������V�i��n,�I=u��<����	�]�'���?Ȱr���땒x7 �`},�|�^#p\�?	�Z8S���P-� ]+���۳��}�;+6�þ5*Y��;z�6[V��pU��{|�s@3ľ��Ｊ׳�LK�P5���̓"X�hE���@<
A	�f���m|��e]�b=�*�ջՈy��꯯3��d����
"*���&է�n�}5+q-���A�YjS��z�]n��Q�N�+��%�k�?O'aly1w��53��~6�r��X^�-��ꗼ"� Cl6=�Y&�ƤX$밤 ����1�փO�O�;���9��(t=�t��ik�[LǭI��{3�e��U��;��g��L64U6Ow�@��X[�Y1+����C�(L.�,{��P���JU9��X��n�_}ܫܕI���FY�	ܝM�Q.z|�l��x�CL���X�������&��j*
���xmూ�>��W�[���*#�@K��5��!������V��^�f�K��_z~�="xn|O˥:vK{tO���H��լ��u���;�ӌ]��Գ���x�?@CU]w�r�x7���E
�l2C�����Q�& g����Vv8,�g�C�~�+5��*�S(f{3�H�C�DǏ$���)�����"�SnضM��i��p<m��>���Vn/�^}�T��+��z�3����P�#�[Kh��y �#�@�a
ɾ�6�O��V��3��;��J�ݏ���#���#H�p�]�(�2�z��%��H�k؍W51"�:T�X��^+���D��\e�T%�4<v ��(i��*�e�
p,(����unY7u5�\���&�YIq�x_-�[��:E��E����i^��@��q��o���[�k���"H�.�A��-�a�Y���#.���۵p���Hם�U¬3������"@3��?�8�9@�L�:�����o��T�]9'T4#����E��5��`wǤ���MRJŦkzWk\/X`���d�o9�T⢳������hm@�|�:�O�5npLm�����: �Mh�q5e�](���LCt�����fj"�/���)/.	���]rf�%�(�*��2
4:�+3�OgEW95#�k��33!��p�����ۚ&�H��3�g�H1wI����&�:૒%�bW�z(�QSF�C��q��v���"���� ֱ��o�����ڣ��Ro���/��V�?���E���G�����l�T(��(��1��X.����c㑙5��=VG������F?Ac���_��u�;z�&k
�V���H|��qs�׎F�+f�~fTQ��	���4�gOe����}�l���p��e3l�i�͑��C	E�;{��5�t���R�!��Nj;n`�^�r�[��w(���/'�/���<C&r��īqWcK-�ѷ#����SwBBL�K9W���6]z^7F�w
�%�?x����?b�@e��P��5C���+�z��O�f����Զ��e���i�G��S9uv�w�/�XΉÈS��F-�5�>C�!�2s�P��E��������J?'oq�9e�EG�咽��vh�$��E�=��AMdbD�Ն��ciz�s����P��S��rΈ����+ވ�Kx6I_U�a���w���D��h;��>V!���}s����#Nj(�/��&H�<�� $�^2�K�f��A�5��3��������6��+�#Ӂ�>'�u�|1?�$}��L�e��z�m��q�B�/�@9z,�0L<2��!�&jwX����Qhw�IK	"��`5�F�c�%EN��L+�j��A|@A������y��lj�_#��(WU2`+"� 5H���Z����J�4�#1S�v�
��Lf�J�8u�/�x���V3S��^9�R��;��'�t�f�T�\X�I��З\�ω��	4b���ˤ�`�:O6�%�v�
l�*���p�G���!����+gn�z��ְ���d1�ģ��ۺ:]v��h�>�+G������c��"2s��$Un���ND��Gf��W�D�?O���tXz���>{���Y0��\�)2z/�^��G�Qsc̥����
���hv��:�h��u5$�*}�>C?�d/�17s�J�	�{�d[AC�>�l�x�2��"�ý`�$~��d��-�����`	��ה���(:�4i:"jX�\�d����ڍ������pɋ(V`#S�K�����~��⽾	H��7F3XJ���S�>���M�Vp�c,zYL%��1��^F�޴t	���s�	�f�����7?���Zi���iC�I�K(�sY�8�[�,�|d)x�\�?���B/�5׽���N\n{��k[ݰD؍W�Uƹ��+����.MX�k�doR�v��,��( RէQJ �I&��� NTe�����'�	uF�cW�+VoqyC�ם�I�K|�/`��(����o�9HfR���T�.'i�!�z��� Ƕ��Iwt�#HB4�ZKtw����eq��"#�O������#�%9�Υ���@�*;�Ȩ�^���;����A2��Ů7#���s���H�v�l�Bp����פ}�@��|W��
|G�@�cm�Le��l-��yz�
����ӫ$��e�or�5"\[�����zF���#��]O��S3�4n]x����7���5E*�����4]ΧP-��s����7ab:��QMy,����)��$�vڳ�VDC6���܊9�kҶX�|`�M���F9�^H�����i4����<ۉR�Y���,�&&�4���7�C��,%W�j��E?�� 6h}�����W��>�w��_��d��-��ɯ����8�M�hs���ꙡ.%�Wu5/l8�/�z��p���,m{��6�0��3����=�.���\�d��&��G�i@���[	�d~����V��=Jh�N�u�pQ����E3Fc�������\��(sj4�%z���;�O춦zg�'��n��G4Ѱw�]�{�5;\���NI�k�葦}3�ExvV\�ʟG�w^��7�Ğl���i=6�`�f�m�q]�_��g�<]Ŭ�fƘ5R�Q�k��v��˲�xH�^��bi4HKN:����'��AH!�\EeF6�@�������C�d���yG������j�-���׮#�����\N��W������R� }fIxL�y�����4�Ħ�`o�C�V7�z�|M��}�>���/��J���g��+}g�껶4�T��V�n�I��y{�!�!e/M�����
�Pөc���H�l-9�{"���W�	X�n��O�I��š/��ʶiS��x�a2j=*q���Ӻ6#��|x�Hx�5��g��y���+��Y�b!�H�Cob����,I'��v�9�s��wF21a*_q���E����=ӏ-�~��
���V6,4�q� ��$�yQ�VFdIGsǫ�-�y���[[埋�%����A��oh�d��~��o��)1�:�>�@I��ZD�as�Q�f�!"=+��a2�i{ϟ�&���e�'E6+Y��_��II<	m�=rIҔ��n^�]��[c����8 &yы*��:>ĵ���w���IJ�e��E�a3-���2���/A-�YBA?�^�x�a����e)��GZ�����{�F6z_��e�q�ɤ���z譞�#qD��D��·�wㆫL�\x���זJ���Ҁ����m�
lcQG+����F����t^!W�v|�cs�Ut�<�"����OŖcQ�ӼV�+��6�0�V��Qw��������m{`�|�)v��\[Yy���|���������}2��r����eL��x��@�0ʼR�o�<�xX��'�%�_��_�"}���=7�#�� �&���b���G����Rb�&��G>.F��N/-ժ˒��%浩{c{��_T���ef��?޸#����ߑ�R�������Q�="M���'Tp�~$V��~�c�hh�ha?|��(��"#4�N���{H�ɸ1˛�����:bh[	b��"�v#��T������+uh����0E�qY%�Yj	9P,ĦH�\������ܹ|����]��ΤM�&@kY��Af���l�ۮKMdJ%Zewq���@ �g߁ �S��
��1c�M}��e�	�7����IL�z3a���C�ƶe���IP����Y�l<"gg�A�o^d�&�����F� ������H�z��QZ�L���"׼f4R�<`D	�l�>m֋J~�0 7҇��|���V�$�m8�2�&�q
"T��}Cy��I���#�`=�e�8��HS.�O�3�dK�;�VC�p�j_���c"O7�,H�U�SKQ�}
~�96�q���\Y�;N��n��)N��l<�������R�"߲ӻ�0W|dQŌ�R���*˻�n�5�1�c�>CfGB6��W�[4�xANֵ����i��\��KN���k�V����H�,���]�vgX�K�9�	S�l��RM�m&���6!��	�t 6�6t��b�=�H|\H1���宮��)ֱnK�[�F��lĄ�`���Y^����Uv�m��T*9�e��t�;� O���>��j�����9��mu�ć��
ȕ�Ay�2qϺ���f���:m}18���{ܼ�8A玲e}��9�gO��?��p�y<���f�~�,P�L�������ɠ�(������M�̺�Τ7=��f'����o7�a�@z�	�~	f��|q�3r}
G��ju�ϼ����/-���b��36<��{9W�P?jv�� $�Ha��_�\g��}�e���'�A�E0��iR
��*�_��`{c� �
zs:�]�y�W����?��'�!�����َm��z��Y������e��Ā�l��4
�[�5E��R�u��y����� �Q�ֿ�wN�S�5#��CT��O �"��&.��a�I��	}״Z �uғ'-���]�W�P����&G����i乨���#��p���h�W�� ��Q�(	�߆�"G0��5���䛕���&`e浪D�cʫd�ͽ��&p<�N��\�W��xp�{���F'82��mWe1V'�LUibi�D�A�+Xa�Ͻ1�S4�r�y��m$5�����(VONk��S�Yq���֛������q��r���[<�4�cOx���@��3e��,e����Ƈ�p��ЮV�3�g��AR��>^@�)!�Å�����X7�I���U�f_v�Ż�, Uj��5'�g�~�d�b�?�N�'H�Y�%�s�Lr-�34^�aD���`E`-X'�A�^�{�˦��'��4��GK�l��-�:Tc�|e�]P9{a�c��Hoo�)�>K#Nx'Gd+�nt�I��'��$!��W�*���NEoysL��.�P�]Ƴ�neR`�Z��ˣ�s�98������8�+j�9_"�+�����84�.Lh�"v>���R��s����x�8���}�N²����c>�|j�/%�=B����G����Po�3|�d�8�%���,m�*���A8����%0X#�����b"����W��>��8�=9�Gr3�J�ĩ�{t�CQ��</�0���p��Lɵ7l81�3@�ҝ�^��f` 1�!��h)�o����p='Ƕ<	��Vrf���ML��Q]/j�6N�O���N�4����iJ��0U>��u��T1�X*Yt�V�����ќch�8�@�*c�pD�%K�%_l�[:+���ٝ�Σ����D(�~�������+w��g�zEn�^��e+��!F��KVQ�v ������k9+vO$����_�O٩z&:^���:س���S���	���q�8��&cgd�H�}����A_�M�2fְ_��N�������f-6�=�^�t��ew�������Oj���XlC+�L%�Л��?�����z!y���s�k�0�@l����JB�!�	+�\�웣mP������e�w��gȨ��������2p�Ĵ^��#�H뾴����$�-F��57� �]u� 'v��zE�6YA��23�{C֘w�O�gz�� ݢ�h,)cq����FQ�PU� ��L�)��ܒ�@(�δ�<�0i�p�F$([V��t��S������2��v�� ��ִ�>Σb�e�(2O"�d������ԸP)(9����j�4^�(6#D�g�'�����@�3���;Ӻ�!BZ��o�OC�~�>Ω��ݫp�f�?K�=��Xfg�]gf��{z�X}N�L1;º��.�+��EOa0A�����Y^�2����,�rf��4�f�ـ%�2��L���8�k;)pқS�!մh{��1R�%2��Ag�9Y��GmrǴQ���{��/٣+��c�s��l��uøDrɸ� Aɟ�r.��rڰ���I|��|���LS|��p���zZ�i��Id%����WZC(z0����M��53�C�g�9� ��6j�P���p;���C#<��O��΄G`^T�'����� 6(�=$�kbF�)d��� p���	 (�,G�Y�ك�5��D��	]z�&C˃)k'��F�.���ׁ&�@�%o��.���3;eSA����f��?-�nL��vA*�д1u��>��
:��3�~C�<@Ӌ+fp��y�NQ�Q��n���BV�@�?�񆴒R|���O�H5T�~�-/z��a^:NBB6�����+X2N5'�U�(�pc|����!ae��R�s�f��[����eqP�hQ�#������v�TN�}e�������0$G`�)--Oq�7�gZZX>��L{�.�����[V�,��n�7�XJ�'
a<
�`VU32|��@��b-��7���>*���
�c3f��H���F���<�����%�}	ϔ�s���� �U��a�}��K��)E�o){{�%�F��P�v1�?q8YУ���1����a5>��VJۜ��b�u�j��p�s��G������=�X'v���s2s̏�+R�M�Y�o����a�����@�T(�G�L#�@�����A���6��M��DN@�g�+�C0dh	�qd��A�!]��O;�m��Q���FW����I�:����.��i��VB���=�����r'i3��655��v5���J�(ꐯE�79V�R����7����VY m�j؜4����hɞ���X�8��6,�zG�g��&*�ϳ��
<�k�T�Y�Dr��fnP+��tګi�O��n���l�0n��Q�'��� �m)��U�l~�h�ٓ����Bk�� 	A��9ʬ]?uE,��lA��G9X!�=+�ى��f.'�%�ׅ�`֑�>`�Jd"B�L+B�t0e3K�JoSaw��i>���2�����(�lT^� a�����d�������B煮+�H: _c��rP�		5��{c+t/�1���`��g����5�^�5��tV��ś����]�ė��5·&�w�{(���tf��P��w-�x�����H�R�Xtg���c]y..�L�v��Mi�� ��8+���D?��~��M�W�44v0�p����Wۑ�m���%�Q-y���=��1�����&�kM� vߖ�J��zkz��֖��狎��a��G[�R����j�/�o��8JI��Ȗ�.;&WToUT��3Q6 ���=�oK��D��hoo0jD��2��/A]�Q��nJ����
��ޚQ�^>��P��~A©��~��� ��p�u����K*�2�q���Q���7��[X���/�"�).siq��f ��D"�����N�h�n7�t.��ǔ1?��fd ��ۺ)��F�~�h\Q���[3�<a��L �;i���X����'r��&�4�=7�,S�5��kܹ9��ԟ��?�"	4��-p7�(��; �9�V�?����{͢~�\>�K9��w����^MGO�?���>;���G����I���	�=�z��@}C��e�����8�p�F�2�������h]��4��%�~s�����T�C�E��Ɣ.�U�3���hKss͛6�jE�E�Yv�-	����Z4g���sW7����/VoZN��#�M�o	[���c��Y����$0��B��Η�P^�4vy�ar�D��W4�sM�:������7�E��Z�;h1z��)�9�C1F@@�����@p]/,q���o��z��4	�������Y<�ڔ3�8���%4Ra�j�ߵ�2/Ӊ���&#�nSba�/�YH�N���^�O��ț"Qgo��]H���sV��5Y��M�FNj�U����"��mbz/r���B�ۣ�(��'q�ZH������ٳ���ـ.�Օ[������/�h]��	�C�rm���	O���Z��
�	�Bf��ؔ�_1֔k݅$�D�ʂ�wv���:Np��+�]�t֖}�p[��MKn4*�N�*�j�W2��~��t�B���{�D<�ȂO?5@�L��?'WmJ$��(S��2PVh��+�����v�\������f��(#����4�y".,x:�0b�þ�,��vpMG��ap� �x:�z����s,zN���l3c�w}Λ������Ǽ� uGQ�B8�9F�r�
����M�3f�m(��t̝O�q��	FCX���l��ӻ[��8GS��};d��Ј���~�^�᥺����7@Ծ��@>ze����g�rdf�r� ��x{d(ھOw)ܸ��l���0u��g �Dw�By�16F8�zrJ�j�瘓͇}n軦���jx>�X#`ԧvD��R��Q�B�0�E�ꋯz�C��۸��O�xU�@>���q�7���E�@�	�-GN�;��>�ˍ0�-�D$��U�a�����=0p0rQ=����%�̃���"�t��%�9��K��<b��=�1B��G��m�ՙ:�p�y�I���}�n��*�k!n���S�E��{{.�	���L��\r4���I6�Րif?���Եw����=���0@K��`��m�m�%�ֿ���7�A;փ�=�m 9QP��D"������l�v�,��jp>]�2�9^�Q�7�Aџ����~���ד��M��)Ȫٷ]�:�&���+�2_7b��f롒�E�"��@�EF!�;���2���Ĕ9���)��1pm�m4����J1w3��k��P���0�y��;��hj��/$;5p���&�c�,o�yAuJ��6�|�*�tJ�ߪ\RKcf���pFǩ�!f�d+*|�!�v���B��r6%�D��I\�
�B,�v�P�0��e'�f��S�Y'b&�qK�}��Hy]��Gf�(i�����	r*� P�뇦�ڼ���a�G\|�gח�=Qŝ��p���D����)��G�z*��&{���	�`���cQ���Krnk�<��|�H��e�=6rU|%�C�W��\�&�����g�/9���%�H�U�i�3XN�x<#FS��:�
��6��0����t�*bR\�ebQ�3�!���AI�ʠ�J�)��R^�0���nؕ����OT�͝����ɖ�o?�|�j#n��g�˒����$�]�\���܃1`vw�;q���G�C����B����!<��t��?	M?D.���ߧ%i偪�SΗR��v���<Dd���ul6��s���Wy�=��]���^N�R�`�����d��s�
Qہ��"Mkc��0�	-%�)���y��e�H ׿�[�����v*�ٞ�4 6^EҠ7���av���:ߣ��K,3����Y'$��p��c�l���qnh����h�+�G���e�w��/�����.�d��3��/��8InP�"��p����6��3��C��s
o]��i�~���ߍ�_9��=f�KȤ�1�����dj�������4�Li��i�~֫L�5�>i��d�3j��0���9g�"8q����Q��~�?�与G8y������y��f��gN^�p�Tg�t�~��<�Y�U�޵���#7��/R�i��U���{rk:=p���p�zpx�\��w?�W�J��$�����3Y>�z�o'�:!C���.�!o�$�C�8t�?^�g.�>�U���'{�J��".�1����3�i�rKR+Sʎ��Rg�?����ߧ�7���7CNM��<��o�\� W�A�2}��7��5���rK��)ĵ`�ȧ�%ȷ>��r&//h�D�-:{�i?
8��nV�J,�mp1���{�x��-�<-�'�Z.ه��Y�EYI*���f�f����2��F9ئ˃:�/ �E�cXum�! �/�C�'�']PI�����[�Vq�s�&j���8ퟏ<�A���H�ێl:G��Q֧y�f����� �|J?+M\>.�K���4r�R��:��m2�k�n6�p�p���4�1�?�]ٳ�ܣ&kGǶ��Wg�Z�_t-�%��d�+N���M��B	���US�?B�URѥ��l�_�|�X2ϖ$M�;���Fx8��aK]5����� B�*)V@O�� [L6�-�bJ�9*B e���&,-?�c{��k�i�m	��.����q:Z��f�Q�Z��Um��}T����Lm���jj�fj5-������D1^��,�χ��7�h��Ω����#m��"��=�/��r���}�@����ynQ?��)�u��S�;���8��(�e�}
�L[F3?}6��|{Nbzi��4Sq�&_�H�-��q�Yܠ?%�����	4ٕ��i��r�G�A�]��2U�N�,��n�����}f�9z��t���|Gʮ���ITР!E�j�/���idb�>ޤ=`b��Pi Z��6��1~ڼE䒚j'Z{I�1鿸�dh-��r�j�T�N�EU�����ր+;ӛ]��E���-c�l#ch��C_��r�����>��M�5Κ�r���$��e%uP(3��s�e��e���F�������Ɨ����TxFr**�˄�P�"��}�w���V�b!UJ��<P���Y)8D(8��9 D�}�5�0���O��wT��i�"�q�Fo|J=0l�9}��z�{��vG��%ҩ6����; 0�� ���I�ݜW���b�?����4��"�M �7�t��2��ZK�C��/����a��?�;���^,JFr��"�|Yߔ��_"��/��ph8]G�#��k3���\����˺���(D��{5'w�(�k磮��g-�м���ع��+�
��x�����'���|�RX�p��#��O6�X޶%xC�����+J��cu�8��ne�)9�� ���U1��.	�1��$,l��s �(��%�C�ȈU����Y%�l����^
�"�t<J��ҮJ�����,YQ�(����[n�~�U8R�Ӓ�'~SAK	�.wJ��kT_� {�O�"����>:+����Kq���_�b=�����se��|������[E)l_%��`�BdN)��:n剭�����Kw�<���;�C�#�c���tSݰ[��]�/���T2�Ы����W^5��1{�Э{��4,pc㻿�U�yN֒��~vt�pK�p�mt����U��V�|v�4�����ie�}w,`@��?���,?�3�b���]�L��nG�����	,��P�/n�J�Ł��1AFoD�np�yP~tpbIK�]dl��瞓�1#��s�V�CL��&B�M�ɫ�d娞PN=��k.�ӻw�!LDc�#�!��n�D,�]h�(�� '"����b�Gq.ëvM��D�N�ȇ��tL��v��5�aN�?����{�a�ԭ��9�����zz	ƿ��Jg�+DRj@r-<.9�:����d��ќ m�?��[�d��.n#c�ŧ��,�C k.@��x��Sl�d��]d�в�c�ؼ����A� ޞd�֮��3 �7�8w��m�i+���\l�!��|H+�%��@K�h���`��wD���%oI��i�u�}~8����V�d���d�s!�_���h|�TW��2�]�.SJΤ���X��[m�y��wy�Z��T�jG���/�c�N��ι�m=r���J�lb{Y��M9K���H.�a�c3~���<���,*7Gϟ�)��q����H�yޒ�z���߉	#�P�����W�-�Vg6�����k�࣭��Շ�/(7N7A@X�u��n�EJ�?k�-X�O���<DL�p����bN^J1����([Ba;e�\z��-L$�����)�B$�UCY�B[-�n1'��"g��ʃ�76	�XBC5�`�'q�PTվ�Pc��x��r�	k�e!�w]�Qt�F�&@Ԏ����H�����ΕT��'X�X�) ��3O���z���	��*_
&k�L�8���%�O��lQX��&Fc�;��#W�C���b�W���V6���_5T�B�
*�A��Ln(�oLⱓ(���\  ���Z)s��e;��$H��?��ʸX@<�q r�m��e�UK���\��u�#}�^wR�a	0N� �2��$g�����f����S�7����1����>�eI��(΀��;���0S���EYȀ�s��|!��^������%�+��� :�k�'G�\3(�Q�_�%')e�b|�ˁ7]^��%еd�̻��7ѸMT���ñ��$÷$U{n���Jr���H��ޥ����<�f
zSE����<3w_Լ����3�6�\FC����Y�bp��x�&�Mg9j�=�����9�#oˡT	^����v��lmz�y�W�֥�dL���.�m�A�x&��Y���ي�t Xh�lP�T�d�cD\�譜&��sjv�S(��?�����F�Hz�s�/�m9?��XC�� ��*^�ˡ��7H-��.h�%���"�>0\	6����'l_`�[@�(��i(�1���˕k{������q�N���?O��s�p����`�=n뢠�p=}���N/���(\$I��;hc߹�
տz%�a���� ���=��P��c�f�s֝���H�( ��# dȀ<T/>Η��`:/cY~�O���#�$��[����x~#��D*��l���Sk�ڮ��u�?*�e�lѻ
��?M�Z�"R�\��x�o�����q��n/����78W�;T���K'۽��h�e����Fb�I���[9��Dz�{th��pN�O�ַ�}rz��ۏI���N!��sCV&m����9���/[��}��ws��P�l"�����>j����"Ř<�JϬ�[=���!�<��B�.?�Y�g}+Y~>�6��{�G�B��G�2�ְ,2j��S2��q��ҫ��O��q�p�ٍ1�Hȃ���ј�����wo�\�I��("r�Dp�ϕ|$����������R��(���	�ʎ!���6g�c&~y,VP����Q�h�=s� �v%�en�oR��g�8��lgR�"D)�hi�{����yr7�<r�P�c��X�3��+�����6C+��4�JR��#����7���9:ft�R����˃�E<ɝl�����,ל��i���VO#��]�@��+��G���۬�@�$r� ���";���:b��R��
�.�@gV�ͮK��ÛId�AR��{�,���&:3��`թ��K��R9�Z58����u3O^s~ہ��
q�G��4J����U��W�2H0l۫�@S���x���d/w���BMx�|�s��a�z�S�3E�^d��Z|�
��;q��l�Ln�Mw��M�e?y,�u?�]�,��vpU����Ļ���@�P@�YZ�L>^�K�\/[7{�_X=FMM��
4�'�m�05M�T��_�4&,�P�6�������-����y �O�	 �'(in�sW�F����{ A;�Eev�t�Y���Nn����q�t�|+z���il<�v�sz P�,eN*%��38���tx߇�c��/P��bB� ����M�+��ʽ���緅��/�Ͷ��[�:����"v�:)�G�#�n�7��Ǥ�}�󢚛BIfB��Ă.���,`�俧���e݃VY���s��t�{ �f����F��[w��L�@݈�2������o '�=�8���8}��4W��`�Ͷd�T�Ж�J�o�9==�#��_@I���)������RWg3ֿpi�?�j��,�.�����>a�2\qu��[S2�b�4�������5oB��F�Ś� !�XqK�p�ڃ���T4u�}�㥻>�}����W\P���J��w@ `�3���d�-�����s!"6��Ko R�>��:g�-��Q]�|�q��ͭ�a�x�-�U��Xy"EQ?�v�.$�2��Ȭ���㤯Fc�V�����z����3v��\Z����bH#%�5��<��H��4O�m@q�r`4KN����h��&ZaQx���v�pI_���yi�w2�]��"3���r��E#A�� �0)V	���%r���(y�'��C����"K��+R��\nx.(�Ci�Ĩ[p�����]P7,Ggk�Xov���a��N��tQs���/���RI_��� �.q���w������������m�&.��U3�d@^m�S;�{�Zm"�xSP
1��q�]1�U��`�cG�X��j��w��o}�&�Eܓ��ՙ1����ř�������ֆp#�>�Mޣax�ņl����q;�<�s�=��Q���&�:R�kot��5�۰��J=�}��_�m��!0�ʒæ�^�Ɵ@�]�%��P5�}ej��ua�n��2j8%=|�����(��F�N_�A�j���'<Q������`5O^�?%��Hd�s��0����A��/���{�scz�1�����P"G��p	��di�,{Ya�_?>�qU�i��Q@-�Ь�[n�ei��\R������Sm:ѝ�/�ӓ���*=�)ǋƞ�����F�z�\oI[lK�OONQ�g�QShE����Z���>�-e{�@�+r��s����CQI>�|�7�Y���-H��\(������>��j��aJ*>�ߤ��,0��ZK�jWԯ���
T�=��5����[R"�ryn֙%�8��Âݾ�9�<�	U]0s3�$�g�"m�W`WA���p���h�B��\:b��8Ny'�������S������*��B�w\	��\d���ɷ�<f�£����L?*F
�<Q�̚��?����Z�g0��?hi���7?߹��mg%�9� ���Z�R���5<�"�32x�	�(���b�-V맵�+����l���t�>ˡÌ�͠~1ЖS,E�
�<~�.vy�����	�R��̺A��g��u3"�[�8����Tt�#��;�;�5��:�&�*/y�[��F�v�*�3�����ז�!(l�T����V�˩rb��NyYr��%Y��}�(f+`Y]�"|��]̟�%�Yh���Vͼ�c�g�Oh�f^���\��Ak ��q�O���"[��
a�|����l2G�;w-ݩ��#�
'�z[Y"~��A���7�d��HB�P�,�e�&)�H�'����Uj?�5�Z�=ʔ-�.�l;�}\	/�wM],�g6��*�CS?)�4�r����_j�N^���f�?���|w0�� �w���p�,�J�����ɮ���r�����:h`Y�+��R��|�)�D��A�bo�1�R1�}�M�ɝ�Y:Tk1�F�C�)J�I��7�p]����9���-rZ�����R�*�0�P�>Bl(6v���U�x(,2��	�K�́]Q�N�4@�{.��9��O)��8A��ቧYCZr(7Z�0���+��W�T�x*w)�]���Ue�Vk��:͊�%��@�(�F��i-�?�s�Ϭ�z@��ʟ�v��p��f� "{��'�s,��Z����[��ٓ=�x�+�[cG�Yü��ep�A8;�pA��*�ca��@�\X��=��KR����#��m�#�{��4Z��n���zA�&�.��	��>�uWo�}(���E��g�5L���8Ƚ���g=�.n-��4�yzm����RV�(n�ʆ9@Z������.=�A���)f����1���;.�Ypb�$�~��^~�����!LX����o��UDP�B�U�<���_d�a�s�.@�h�!f���H]Ǉ���H�{;E�W佪�-�4�O�.m����@�"v�{<���E�k�Mv��x;Q2�>E�c�A��=e��$x��A���,4�楓7:��k�)f�C��j�����"}����=ʨ�sy��=��RD�r�zS]��wPw��n��F��ō(ݕ��Uu���f�t0Dbs_�JGR�*� �3�V�&��F'������lf0<FE�MQͶ�ݠ(�*���/2��)-��hg��A�<�4��`xf.�mS-��,my.*�s]���9�E .��'��,R��F/�Q_?X�B�L<zԍP�y#V�LE6�����r��6\٧?��nkHR8��#�C�?�)�yfN��=�u�;�J�r@"�p���
�2 �/�yJ��*�b��݈�E����lm���<� ��&�'��Vc�YF��ى�k�Uל�����ك�4��yV�n��)!ͣ=q�a�0#׹OgK�r����dV*��L)t�'V� }�E�%�ϱ �����z-��z�a�
�%f̗���j|X��,��ʴg��Y�P͟^�2��;��"!'��ğ�*s#eg=��^A�GoYd��o.��к�ݪj�a��ã���k��\���=�GŻW�\��nHT���ee%��l*ΐ�},��^��K\���XΫ�q�EMN2����[��p޻�ahm3P`}�?,0n���Ї;�+�cH��N��c�E�Duw#5mD$�t�˞9�ڣG;��t`o�x8)e����զ޴��{�ϸF��c����Q��[ �����6t������ɢ$��yM�t)�T��%���r u��F%;���P�6H�~�IJ�w������rX6�����09r�s@�+B�`6d�	�����I쾆v=��V�YP�p��/��p����Ԯ����X��!������lЩYr윳�ы{z����,s�4X��Y�jcPu�A^��r��ԉ�퍂Z�����_]�}�QՊ��Q~yGƱ(c(^��!�js����i�,Maj����> �c���D[���OU�%A�s	X-�a��آ�b=��4�9�I��׻��1�����XO"���#z���NK��*?���D�p�����Bޛ�����bo�!4M\���-����,4yD��">�:t�<�}�������2��!0=��j|�n�o��Nz��-޼�Z�ToqG]�!���Ih{/�`�6!��Y~��>Vw�K�u!�ltar�����4���QFa� �EM�/�d+��-����#�ɇM��\BSa��O�W7�4P��N�o�ז���uF��x5�K����?$���q���Z��xp#��`���?hM��O ԒD�#�À��(�����+�K�ђ�!s���UC�gm������;���-�l
3���u�l�F�ᔈ����wNY������È!v��q��>��W�>3R��i�Ι�3d
�;��G�)D��VևȤk�ט4�ox��>�8���՛�8�jb�j˭�_��'��n5qT�t���JO��+yu���0����y?d���Rs�˖؂�34<`��7�«)1㽟{�g���)睁�����^s{�;@��h
�޾�_�?�Ј��$�tKSFɐt)GNhsDj2�0�j�_��0�;gJ�yHĦ�gH�Z�}s�����
����n�Bƕ��O;f,�F�AF�nH� 2+5A�c�@�Fv�����W��G�E�S� )E��m����vY�ǓN�L�肠�:�E��2S&������	T|���#�l��K��A��Q}h����V�F�'~< ��0�x�w�$�#�Ť��9mϴ����)r��^�s�ӄZqm�vfǤ��I�s2�0pf65�`=���s�<��{��!�^F����S�@�5901�l��>3�}P 1����'p�ó�	�º/�+��s�p�xk���ox�ƺ���#�}�"�U�H�u��W������ �;�d����rЃi9wS[�/�9�wbY��J"��p�%�3�Pq�,�	bB5���uӦ½g��`O3kٕ�^p7���I�X��I�H%GW���%`6���q'��&$���WfA����˔��n	L4Ը������.7έVnBd�yr8�x�g��.�H��s�WP�߿3�o@�[`��7^du�>N��۫(���6�W�q��6pxX��N:���X�)����� ���g\��W��Ql]d�uf���6�ܽsf�Z��k�QF�n��s�Y�3h$�7*�_mQMl�`�+��N*���@�gوN��6�ͮ�f�yOd�������8���hiS��<b��kN�b3_���-Y�)�d��vp(�����c�ȗ>ݸ���KԌf=�5��J侶���p�y!��Ja&(��a$���L�.
������Sc1+�7��%s1(Mh{0+�-�w�i�b�A仛���9��-��܇uk��By�xTW_m�a��%�=|���-ƚ�>ӏ-p���mɰ�8����c�`�
�iI��B���;���pHf闏j0_�&��}<�o����jG����Ta�m�ʸ|N�x����TU��Ѯӌξ+ęV�qo��hΪ�I,LF���B&|#��C������0U^�N��x���C��? r�Լ��h�O�$?���q��֛5��e�L�=2}� 8���ۯ�=�3=^1�*�/%�(s�9�J\{��ׇRzW�R��������*��N����x���v�	(�0c-R��%УF�D��;��>ˇ�.!MO ELEʔ�ȱ�fd�1�E�*����iS����:���L�YT08��T
�q$����o`�7p\��`�܂B�z�/�Y���r����p\9�{�k�W<d�H����v&�6�V��O������c�<�3Q)U4J�rD`w��󤍚4���	?~5s�%1.RG-���8�`�)�'�^6%|�[+��j��r���,"��>��^�Y`��>ȇ��B���WӤ��1[�c`d���?!�di�'��e�p�7Rԛ�\	��!����ȳ6I�Fg�@PX+K$��}:�檔��	����08��)��,9���'����Qo��ȾM9\���|���m��"�po>e�� R��x��ѻ�ah@D��#���Hf`3��W�2g�-6ɺ W��2y�}&�5 ��'��O���7�m��M��÷q�w�(���|����@�G6��U�:i3p��05�#��D�ݮ%�Oa䨒_������;�Kr�7�ܩ���s���9�X��۸okT�/T��-�i���K�\��wn��x��F/2�>.�6]�(3���+"A։B5N�1{�n�S�&��A��[���/L��p���21�?5-�8�¦��˺`8CNሡP"1J1-�m&D�ң�Z���R�L�/F��2r��0_(�&�����{��iƢ
���m�Z��p+و���y�]�U�0N,���Z�6!F�K�j;lr�����Hh:=��6튢����p�x�=���QE�2���^�*oᴥ�6��F~9��H�K�Za3z�ϸ�}�e?��Yv���@�A��I��2�m=��`�0'BkTט�:)�4�z�1<�|39�O�=�X�r�ޟBO�̛{�\-N妢��tl !u���D�YV�j��B~�I�d�wʳ�`=ޣ(�1��^����� ̼Э ����WE��en����)��Q��K�׷�ɨ5�Am���Hw��#����h
ҏ���R��w��]SoZe��N��섂��f��s�����uRٹU�4t{�#5$O�n[�'GX�02zvЧ��Ti5�@�d��u�M�32�ܷ)���VHa�)lw_�+�P}�چ��H��˲O-@�g*[�� �7��`1M��{�3]�X�E\/���:^�*��&�����'Tc����������O���}��ʴ��hW�Ən����/��Ez?��"��-���agO��Q��m�����&-Qȹ]Q��oC|GU�)G����,��S�X<R����@������[��I<�^���K[$v�s[xF�[g;Q*�\=�"-��;��ٶL������v���G9�k�3y�-���:J�r���T�Eh���4&�`)�#�,����7���O�,a��`u� �c�0=��	�aTg钏s�h�{����#A�ZW�� ��;�N�!�ED�ڿ��
Tý�w���4��o��]r�IX�
e���9T��H�k=�>o���n�g����nnA�ml�nJ=ĿM\V6�m��	��4.�#
*���h"3�ض��9$�)܏�˻���.N$�N0�X
��N.�J�`�.wɔ���eJ���)��6��N���s�=�`�9|K$z���7�_���W�^���P���8 ӓ�%�-<��\'�,I
�(�$0����%`�l�kCV,�u	��V�	�B�{.�˅i��
�d��\�mE	%�L>ڸ/�.�k]CWi���Ѥ2kCZ{�����i^�h:ɔ�T��Җ�����Jsb��w�B'�:��4������W��u�G������U����7{Z��0�	2v�݀A�@�7��KZ�I���̟"�C�"�tݨߋjd(|����Uw��� ���z��X ����ۑ�!���9RS���0�/i��ȱ�N�-@~�-T��辑����"���D\O���S Q��'�<*`�1r�����Zuz�Ƈ��|
������EW�&�B�"�Dj�)m�R��Mm��@7�IKVk�[]`�Z�����\n��oб�&�%�h̼�����p!�	�>n���qa���q�I$��d����uQ�@�LiK=���vcP�����Nu�~��l�~ʽ�\c�H��W�g2ь!���Q�-5g��ҰQ.������A�\\�u}�� =��K�R���(<�D�Ɵ�&t�q���TM����*O�'���N��j�������,7���y&��I�"C�1��P���&e.��x��M�|."������g���4ξA֜]8=W�Og��v<w�ygN{�yg��`:�!��堕ev�7
!���ebz٫^{����Sz$/>o��N�.��d-(��v3t*+��Ղ��]@FAZ�Ң�=Rh���E�Yt�`X� ��b���@o�k�N�/�@Ys�8�!���B��LĢ2(�.�O�è��'Fe'�N*����/�\�^�8��Qݾ䟝���:���|%m�V�<�+��ax����1I��;R�KD���$Mqk9[r��÷�#�aVg#����m�~}�[�iq��3���E;������$����{
�{Tߟ�Pi��lt��9
o�I�@�݂�Һ[_��A75Q���CNJǹim�� %�	��0��u�S�P���>�b���!+�x������W1vR��=5�S6�yP����k~Wѕ��8�˥+��o`QU7���^�h�*p�Mo���ı��H��Xܖ����˭�!)��`de,N�П�J}��I4b��E�̯���g�-s��|�
�"[vV!���~��6f#~���U��P��� K~�{u�s�h�j�"a��_?i8���������!)l�3#�P�۵<CA��袿�Չ�c����ɗ�I?ܬdR�On�~����26�6�A8؟�Le���f@$/�C���J_ǃ(�����²�FǏ��1J����� "HS5Dnϸ��c��kJ�1����*��SMYl����+�<��2�>T_�_��EnF%�F��`��� >.��9��<�C��n!;��.��^��u6z$]z�>j�ᐯ�cc����'�jq=�b����fTb/\�xa:&"H�!��j�ۓ �V�F�P5,��ͥu�`MT#��p7��t��!���/bv&jL�G򳕵��oj4��Ǵ|	��M�.泶yD�"ci�|��[A�ڸ,�������z�pcq�\e�1��YB�P_3v����Lķ�yoqWTj���,Dn�0�L�B�щ�{�tZ_��_�2�����y$�l¨7�J(�.�E�����_��i�TF�U���g�8~�<^�;��U�L�4�d�C*;�0u�1����x���쑟5�X��-����ͽ����.��!�W�^�v��������U�:�,���܊|X�����l#��(w�ޖc�p���9���}ttG���F�G�g+��Rhxw�M�qhf�?7���(�r�f$A��h�&ND���پ�oPrRJ���K��x�M��)��.�e��� �w�aMd����˭2vܪ+_��M��#�ӿ_�^#�P���Q/� �"V�v#��U�L��=�x�;Y0r9`]	���B����� t#W�5�w�⍓Q�f�\L����_�_�����BE�ӕ�kf2+ٱ��F�����+�4h��eSM-�"y����.h�O(�� �M�G���t.)5�}ڃn1C�P:����wU���1{��*���8��K-`���V0��5T��8�i���z���&�y�夦���v���P����G���j��ɝ��aqJ����찕�2�����D�Z�Q�l���)����L)���I"ys]�)#���#�����>�6�]Y��8\�X��5��7�YTg�,��<���,Z-����gv��Ȫ��RW��vFG��鵬ߝ�}ogn�ES �g��i)���bUL:�f������R�{<R*6�4-g雑t��mv6־�e)|�X�6�U�ȁ�M��T�ޜ�#�bA�
�ŵGPS� e��-X��T$�����81��v5��i��M�v9{�3s�j0x-�"��\?/09].��y�� �jOP��r��q�-8Y��8̇�y���Nj@�_q����+0�dt�0���0��������S:��4��$"���g��˲�������	�����Sz��6��hK���c��ۊg<��� �[7�l�DIη��l�~l��?�������;�&�C��㭝W��Aq�q<�ÇG������zH!P��6��h�Q<J��\У[�=@`��r���\]�ˇ��\Pa6S8���ll���Ml�Td�
V�2�k�Lf�e���~7QC�K�k�$�Aq�rl@��X�۟����/ �c)����zKÒ�S@ń��m��rݴ/��D��ÀU�]��ma�(�ٰo�F�W�ia��%|M g�*l�b��E=C����4�CPj@�)@F��;���,K\����K9z�4�V�!����n��U�fn%��"!�L��WΛ�+��2�2�(z<�hl��0f���V�ל�[��Zd�e���	W���l�,99�� ��#ME���r��u�e�\�r����bU��TKP����!���T��K�"�������8�MV<��H#)����=v��E׶E���ևp%�[������a";P���N�H(}�$�,% z��b�{K��� e����l����wK����:�����b�>�*j1U%��I�喷$屳8w���R�8[�����*](rK�&(�Q��xe���Vl�sl���K�\�I{J��,�+�8���>�徵�wF�D[�XF��q�`��_��c��keZ>�=ߔ�n��d��N}W�g���"�`��!5�7�<��w���kܦ��� ��H�������b�$u���k�!�D]ב`��xx]�c�vZ|��$�z)�q�|�B�'pB�4���8D���A�p��	�vH�k��=��I�e��SK�G }�U�	�*\�x�k�̪hmo���x������f���Ú��Q+i�T�!�W`t�����+�t�F7�T+�����heG�X?����X���}��� �'�*�О�A�OO��4�b�P/�爳Nc��~�DC%G&��3���*��g�#X��-�x��rJ�>z��- ��	��d¥o�頻3�d�P�=��/Ê��v�������82��-MW*��k>��Xuh�~f�;pA4~�[���"��Q��1){yt�x5��S'�ou7��C0�\�)��\+�y���*:� 4���h��o�3HU��q��Oc����4�Kd���k؟�̳�k-�'%�,nU.�� :��G��wX!���ȡ),_�^�������(�
��)*u�
A��K�՘��P1�Qq����ᐟ���QG��X��1���2NYS?��{���e�#�:�e('��X8�V����F�?� �3�r�ŝ7�a8�V�,�I�]K�r8ޫe�_w�"7�d��`�J���L�js~��j���(IQ@�`Ѷv���me����~Z��x�h�.��S7�)��~;&�6���ʣ.��#�2�k%�m�H\���'�r:�!��aI�z%��l�:�� O�<��4h1��� ��u{�ka���<��Sڃ���ߠҋ����96������fz���z\V�Q�R�(k~j���� 0�Q��T�����a햺:�l(���l4�[��OP���w`���Le53S�o���%�/Q	��-*��x�W��R}���z����n�8*��u�R� ��$�aY�4�$.i���uְ�'��Ոv�[5|�*�J�B`�M	�c�f?��2"άM]�n��q�@�G=6�G�L��ȩGl��i���h�z���x#���r���X���/�]�H\H�zOǯ�W���\_�ʛ���s�:�U3	S9�Zn�K�'��Ց���>�x^e��ī�����퇨���[5�Bz�1QQ����OxǈnY��c�h�LM�J�a��Uj]N����*0|ؐ���\�R'�hAY�dz�Dr�V��@�8�X�l�^���#8~�A���"��\W��WtH���G�/1)�}��ֹ�z����S���c=��[/w2$nk��K�0b����.�w!�y�f[�iڻ���q9���4����8E��r���+��I0@��ig7/O��������p����(q��P��*��0��}��k-����Ͷ0�
z��F�7��F���U�^>
h��@�������o?��� P�OC��Z�����%j-���{�����p(��[�X�F����@k��]jxv�	���?�~�<��#`9��(��r_ED9�2{
��!&Xf,�I�{���� J�E���߸���II=5�s���1$i���%/�#M04Ar�͘[� =h��E�1T� ��^q�є�9���m���=�hB�E�9���5�������G�K�=��!bm�Fr����T�Ȁh�҄[acq鰸Ð����x�������]�54�ܔ�U[��"?$����c�F/��v�_I$#��ңZ$�o�ϝ�G=z}�����E��Bh�bu}�[N�L��K����V��4속lu���~��޶:\Q�ۀ��m	��l�F߶��������ZX=M�>+��l|.E��@]���A/�5�p�ls��i;7
�G����~I��언݆Z�;x>z�M4��ҝ�V��&�'d��_������QW�D�tA�3�oc ����fهe��r��~��^!xv��
�uU�H�4�~r�xq���6�2+�.���q}m՚�:��+8���T"l�tf x���#;Xm�Ϡ8��UդH�=���xv�˂f�r��j�@jԿJ��8�!�9��H���i�{l����{���vpl��A�6Pܰ"Uy#>�������5[�h��;����*`��/R^y�[�y]�lBi~J�u(�M���WtO��?��l��6�ɐ���[�R4���I9$= )6�Ms�F�j9�1�d����mq�p�V�ICS�L����Ȯ�n��������6�P�W��:ʓ3"]�ɞ9�]u ��g��I޺��'�y ��;�/�����r�,�Ф�Qu�]�gC��s`��~Id���Ž���&��\��l2<^-'�s���SO3���N��.��.�{+5f^��	�3ᔏ m<'�[s�� ��ig�\�4Rxd�k��Dϗ��ޛ{OF5�BNP�W�8� -�3�57g	��` �&��H�輬O_���w�P���~0Y˼G��k�g�vc�[��Ɯ����m(�H�u��Y�q%�Ûl^�b�x	����!�ݧǚ����-:A�a 竒�����c>��g�+t�̬��)<x#������_�S�p)ٌf-�(������SDfC�PC[IJ�LΚ�v�����Hꘪbe	�L\�au���� �ֆ%��(���e$w���|�ʎ/Xq����s�y!��fX3�[���5^���i��^�jc"��ˀ"����Јy��$zQ��hf��B}�  aI�¡s���cW�P�zhQ�WΕe��Er38�g� ���L���2�p��U+�[�%��R�AQ$�]+!W�G_��,l�q�����L; �n�f}!�i�g��3╔Kn�{���j�D�r� V՞�б=��B�(��!D����a��2�~�~��U��ZPB?�b܈�������J��?�h�W��=��;����"�5��̐f����ή��3��ye�ʺ�����d�S�;3?���A�e9v�#����d��~e�g��	�i	��bӗ_xc��)���3^�T中�,��zl�\�ل���{N|S�p��m��d����g�C��3c"�@���b] �"����SEB .���Z~���>�'f�Q�(%'�A;Y\�Jڽ���Ƹ�_��_Lٌ-!ǲ�����w�c�d��*㒫�E�|k�h�瀭,�
a/ 31�;%9�47�E&��W��[�1u����p�~Z�9��C���OPl��H��Y1�,RЌ=���[-�ŭ�?�o��b&9�0�}�`k���2�8*��s��˻l����B8�H���Z��-�P�ODb�؇��t���HZ
���y�{3D�LY�GW�	�M���kEr�z.j�NW�Q%˅�����<� ���a�X���	O7!_0��re���tR��d8��*��� �����&y8�>���`���0f<������ �ER�LC���^f����g����X{��?�	O]6g�+35��A���
z}̝޹�!���p� �ն���sp�w�|� _���F�@N�p�V���f/��B3|+��S�vDa�p���8����ف�"M�����UE6ksMsG!s�݂ մ�c �d��!�)@{��S@�&���v��
��n��<v�Ͼ�z��.Dl!>��SF��7p���q��F�!�����������V�W�ٷ����&DbB-��zM�Q���\+,V@v`�.8���Y)�o�.M�K9l_4�ls6��t���B�E�j7�f�4dn�F���ѓ����� �1I"���_'����)�(��T��Q���l����_��˖�'|�����H��2�H�������3ӍQ������c�1�h�W�uDC�C�R``�G	�Ά
U%�>tJ*��˒Ap�V�dmsB|x���VKpE�� q��w�������]l��i���	�+Ĵ��]4�AW�R�eY�jG������@<��W��]�`�\����]W�k��6/��p��aC�1�[�N���/>'�E:j��Ȇ�a,G�xZr�d�9��A�#}�@xז�h�H�HC�h�H��k��/I"������,�)�����.�m��a%��MC���,s����x�����w`�����r7R�(�J�м¤��25l��Q-�����]���.+����WM?�3y_��w\獷�炣	@�c�G`X<�Ҁh��ϪA�
6�Ѓ�-T��(Ͷ��ٛ;Z  {є�I�*�IG���ơXo��⸓�N#ޮ�)2t��+G���߆I+-ݴ{��yp��l��j�q�&]��=�b���i_�����v�7>~/ƫ6���e��Z;���@�j� o{?���� K���>�q<x��1�H^%[�t�uE�Gx���u�%�w��`����Q:���ck�k�r���-4��b���k���e�	��C¢^*�>��~2HA{JFs�Y��v%��H�챝���/3���J[�W9A�!��|�GݵY�)�~%�<d	�7�ʑ3X��ǽL&�V�+?�w��9o��@|��3��1�g=	/j���Z�[��(Q!~ڔ@)�e�9T�3�f�0!l.ًc�6�9Dp����2Rq�}ޮ��wJ>0��E7�aIY��e*�	k��<�2���g��g�N[�M�k]\��z�Bv/v�����ix��ɡZ��c�o6����Z�rS�{)81N�@ +ͭ��nm��b~ZwO(�iH�+��^���vg1w��~]!��V�5���)a�֞�Ќ�<Jr��A5�(��"tb�k���q�lWV}F%N9̎N�ۼ&���`�V�f�L�Ҙ:\|>��G���2��5)�f�(iŎ߃-T:�ZvFFܳ`����;3��:Ϙ�2��m������f
!HL�[y ��搒��u�%���͜F4L�b�yb(����u�6y�Z�O�����;EI/���X`Q���D����nZ)���������'"��r��fS�R`��H���.Ŏ̬	-���0�.Yʼ��K��[�.�Ũ\x�Ft	4%��oB3�$1��`ǯ��9��wl�)��>w9vؚ��z�f�{�;����x�G�����1�o(�ʩP�% ��6z��a%od��!��c�������=IB�~�<;��?C�}&�����C��zSB
�N �!�j���&U��Q	�@yw��
����ܖ̛���֓L�y�8H5��̢�z4������!�-}]�4p�j��BtxO�4���@ՠ�
�"j��o�}���z;�ii���} <L�2��T�z�����D��D�d匑��y��;��D�q��<1v��"c7;�]�UH[d��m�5��t��rN[(���e��aOD����T�Kn�feA �\w�`|�rt ݽ=��$�g� ��"�w�����RԬ����>�:k$������|&H��>�Bp�W�S�"SA����/-�<�O^����)/;��o��Y�(l�Ps}�|���l��:����ߠ.~Y���Dz�ew%�=ɳ���5�3|�Ɯ�SLʒ�ԟ���o1���tp�2�B�OD؃)C��:bD�%؈�����Ґ+��tV�ԏ��'����[��~�S5�m��V���v�%�j:R��C��rz��C�j�A�{�6�ݱ]���dcl�C���P����;�w,�����>إ���H2���/��Pwq�{i��oy�ɓ��M��f�G{5��>�ϋY���#,��~�L���x�S*�6u	a4��q����f�;q�Fa.�<B��������E����Ò������L�*N�H��S�m/��s��Gh[![6x!�C)�[x��{k��|�/*�5���~�Ke�<���+��up].�� ����N���?F�`U�B�"ws���b�'���}��m�٩9���?!!a�Z�|ct��G_6��Iq�@n���(0�Q�#��	�� �7�Fb�a��8Z��ei���?n�|n#���X���Z��g��$���|��md�A��3�W���<e�l1]1I;��v��]7����\�;�,��!�	��1�����(^�9�^����/���W֣��Vu)��bj�9�]'_��
7@��6��X�LZD�t�wa9%�_v�� ~U��ӕ�K�_d�S,���iH��u�w�5�@b-���e�0cu_ko�iK�3���fZ��p$�Hu=�6��[s����0@�П�oe.t��)��Ip���&0H��!����Vfo�Տ�b�S,_�"n?T�힢+(8i˩-�n���^S,�!��p��Qḿ��TO_�J��!Q�OM�ӌV��s2|Ih���O$������k�J�,����p\�C�"r~*]�jVeܿ׎a�7E֕b��n��a�q]֕! -�E�����9�����L���M��M���E���h��:��Tg\E�d�i�5?���;�ҽ��*6o��T�&�=
���?���F�cn���e��M����6��<&q�Q���U�y��U�f�;����v+Z<4E��J���#м�u�м>����8��3<&��}��Hid��Ρw>��i����o�e�^��;��?�1�)jQcQ>pɉ� aX�Z�� ��T�V� T�ad���.�4ɷt]-��IG*���s�&#��r�㼨ԯ���8�[�ڱfg��@�d�~=.������y���OL���L�ZDYyo�@��(����å*�4���޾?�u��h�)Œ�L$�!6å[e���OS�	��H�e�,�,M��0��^�K��+k�F�Vit��RJ��jU�)E'?�VCs@������J}�^�� Wt�"��3�j�H���C��d�Z)}�2��`F����ݢ�Ӛ���2��nAҵ��Y�{�g��TK���N:'K������~'x��\Cܴ=��.���$�g�C3?�V��-�V�V����Q.*�Mc�J:�\���E�M��@O�ndS�߫6ģ���D���b5�d5c�a�mY �E-c[�+�u��u��0NL�oޢ�PCI�?.�����$��Tր�؁�|�f��׫z��T&��R�3��.�SʿD^���9��$�J���]}��9�z�J3�y�:�=�V.�	�J���HȏŷԈɂ��)����
wnHQ���2�b��Cݿ�]6��Tf�F�Hl�?T%X�ߋ�7{78(w`ɡx�!�6M�+�.��"���0֐0À�F��+mbS+���=��#�`��8=~�? W{�6�꧿U���P&�B��3�°Z
��`rF�H���Ob�CJg��`-�K� ��p�cC�_t�ݯ�Ze�z�R�8!�9��/�
s���Z���p�O]��*X0id&V�����vh���˻�C�l�?�V2��M� ���稘��m���2wغ�c9ʣ��d8fd����Wm�"��@�5.�J�<���R�Ff������ �y:�kfۣ�ߍ`?<�o�=."
L��q;�ɡ�!_���f�-XL�,(3��}���G ǆ�w�.�P T�δtZ�W�B�!ܑ�c�U�ߚu�z�Z�qqIE�s���C0���H�3�bK*�7��,��p$�8i������KD?&M��9$&�PѳB<�����brI'@�`0��NU��.aF�&]�t�Cwr5�l�9�I3�T' ��3 +�CǎZB�Щ����%���
�2`��U^-E�����C�T~�ўw~ឝUj��u�����1k/,i��2�^(�u�I%����TP��]����ߠ�V�'�/������b?����pz��]��y����cO���hˍ�JhrnCg������V� ),��\+r�����3�������du��<ԥu,��t�]+�j�}�3Z�����~H5<���|�/.�v����h����R��A�@����;ʧ^���ѝ����lkle]P p,8�^�_w���5<����^��U �k-�,�6��'�%j����ïIf�ZBa9'<����E��ZJ�r��X�7�A�3&�E�)`p���{����l�͵��M`���U�Xb|x':�0�����`��,SC����H#s~�����_ʜ�{]�l�"UL� h�XFJV�j��-���P�g�rA�cZ	�ޣ��@�k&mb�ҹ������C�pǰ�dc�j�mt�2��O�8΀چ" �>����͙�� g��p�Y�}Rv�V�&�'�cE�V_�z�G8O�.O�C/�Y.y%1=Rq5�;�a��rGjyK���*x�d��&9����m���,9�&4x����;ʜI���&d�5�f��3��"Jj� L[���^�Ղ�]��F��hH�袌D���QyԲ_a���M��N9����f�
R֡�.�-}(�/��W�P���������XW��Q����yҬ��?>z`<�9��h��<-p�P�a�8�DX� g?Ҽ�J�n��D��'����̖d�hMu��t����V�W Re��jXk�Esݡ�z5�*�%����z���b��kS�j��F�
F�6;��<��f~K�g���N�g�]�}?�W\�N����)�ty�Y�����1���W�p���2�/F��H����*��$�ч�p�(�����S�o������y8:�eVL�����,��=��%"ű�I1��6Ӄ��ZR��;#c.��:ڥy�M��������ǧ/u)3�Q�V�Ć����N&�΍lB	�f7j<��n5"��G��It�i���4`l��P�AQh�3>=o��sn��wz^H1JE��z�շ�pR����jf�2<�b�.�Pu��s�U�"�Qa�p#D��*K��H�F��m�D���\�7�V��R�i�O�໏������ϋD�czE5P��� �ZT�hu�̵��m�$B���������*��a�3��[�7ęe�H�b�:��G�'�%'��sv�����w�`��a��Y�ys�m|��,-��������Bb��	���
����ǍO��|��fߙ��ɂ���
���7x�G����G䜭9�����;��Ω���}{��b �G��Jo��#�<��DYL(�=�
�/8y�BD\�HHV�bƙk��xzXoY�������B*՞�ªT7](��gbVѝ��Sj��٪9�B#U!(.�ܕO8S7Op/#u��3!5<��1�fߝ8`
����
L���Q}�6� ��O��j�L���e��%g&���f�� �a�(�O�)���DB{��H�L#{�)<����)��m�)������`M�һ�5���S8���#��i�7i/{�t�Mӫl�5-k��� O/�;w`c�wxٍ�t�Ot�J�mtN(�=��/h�0�Q#S��x'�h����v�\6o��:zy�>��d|��f�	��g�E��[�a�&J���
d�)K?����7/Fy����W@���I�]�SV�Ai�n��8�L�T}3�v���1�IҪt�u�~J�)<G^Ov���i��W��RR59��q^��Cv���rj`b2�W'K�k4�t^�O���`S:�J��vl��6���@ �|�k i�������J�;���n8@�HA-�nJB���"0~�!.Ј�D��|M��D3+=��h����#S:��ҹi�A��[�����=���v���l��6lF�G��k-C����S�߈�Ck�7
��d���
�lP���>phSh$��ϝ��?B�5y��qO�#i�a~�h�s#r���� e�V�9��-L��q�����$|S_�b��(P��X [��9���F`���K75�mh��V\���BA�D���u�qw�D1�U׬$s��@z8��;���9@Z�s�A�%^��?=6v�����ps;֠�J�ۚ�ܥ�"�+��cY\/.��3�p9c�	S"髁z��7j���r�"�FlU�1*�*�1Aiu�1��Q����g���>T&�D����Z��7�{I�F\��{�x��̇Q��~N��v�xf��|��xxΛ4}݃WX�l�+hR�p�P�1SS��RحJ���!5֢&��R(z;�9[˙�\6���[_�Y>|8ԡn!d_�جeY�������>���Q���Grx� �v�z� Un�J- �� *$��R��ÿS�E�#g{pcA$.�u�%��.� ��6�P	���eh��>�ۢgw�7�h���>I�W�3`�WшEO���FG�ܼ�ˏhc����"��Lё��gSq�����6>T��1���E�;S�x�|����>C�9n�h4���=W��J��$�A+�0���=����K���a벪����o�FhZ ��*�Q�(Hݸر8�޻8��n��^�����5����rȗ'�hJW1/'�=��0ܰf�ܙ��N�]�ѦZ)��U�vB��i���;�N�?����e���ʰ�ģ�[�>^
I���U1f�^�#�([B-���gE5a�f�1� 	9A��r��]�KT1=�%��i����_�7�M,P2'Wu���Q��;�.��
KX��U�]�+�Y}���.j����P;5l=M����wK_�aB���#H���3��L9�������#�Y�T��2|ypt]z�
6>���UU��7T��+�$��*�������z�d��kE�(�Fa)6j��W4�)�.��VW W��%M����x��!�D�UkVw��۾^��O42�|C5}�F�j�-��s�y�M���g�N���w#�W�m�l��f��h�-b���:�&l��u��n��Tz��ܧ���/(��+��}|RQ4Z��ԏU(�z�Tm�<���?��8=!���\)��ކP��jy5�,��E��J߹R�a��Z�[�xg{��a��`ŪI�JP�\<9;~�[~�� �h��0��p:���2am�/���28 �
�{hw1L{�c=�h�z,���Bb�"�}�N��	o��x��dh�	\�FezΙ� �,�]n�uѐ�4j�^�B�䎱H�G+\�� UY���ID��� X!:���%-��F�sc�d/(������C��+���-��L�}���J�U3oud��@~��p�D������p��j�<J���f�	�3�3���=��E�'m|o7�@����?�#/�tX�3��l�XF��D[��F7ETj�/�'_~�KS���Yn�UWT��
&���ӆdo�@��<c�^�O���ӓ��N��C���z�~rKZ���+��H[�j�� UP>���]"�����(E��d'�h���['��K�2�ay>-?:+L���ުܚQ\#�r�$�-Nuy�)��=�!�j�8s��U2��h�Ǚ������t��j3&�u��}:y��l'z�͓�⺑=��?:R�>D$�����	��;Q��>5��}��|N+�yW,�w6ۗ�����^5s-�PO��U�D�)�}��\R�Ghя���9��B'����	�0��7�4�fY50�,�\�ͦ�C��H�LL�l�hq�S�#��Hi:��ra]��wF6�~ؗ��S���F��J+��w0�Kb�*�����N�8���`)z	�k�h�9��u����ADm`p�d�!�QqB��*��U��-'�TM��8�a0��m����R�7��Mǎ����AU`���h.'-E�3f�LƸR���Q辸41��7- /�
u�s̨��4��,�� ��>�]56j�pʞ�� �}�n&M�.�}c<�HJ2�������f�IRAI^�`��N&6��(���o�"[���,��җ�o�u~ f�@e��c#+�#���t��$����!�9�rL�f����	��M��!��ӳ�^b��[Juo1�v���*�� 0��3�%2�ݝ3f5�}��+m���rB'����^��b�э�ze���DХ0#N�`�F�,�u�ļaRD�����WE�d(=��P�sB<pf5�h�����g�C��Ā1M�\��z��%�?��ʸ�����9��4�p�|OWȈok%���d�u������ު���.����p�G���d4�@�9c3	<�[�~W�$���X�Ԍ���ɷ��N��I�^���"��3M]4�%Ʒ.
�h��B�Mf
��������Ğ𻢇��s���0'��t������b�:I�Ge�L��������o�=�  &���G0�т��u���C&�����!��J��R	�1(W�s`;1C�;x0p�pP�z�o\k��ll�l���]'{�2!Ed��1�X���3!}�.w�֌��Yj}ܱ��6���w�'w�z))nC�r�i¡C������N���1���­G+��?�5=y�c������ᡜjM�U�iƯ��9��13�N��4}����3[�O�?����N�А�^�؁��x� �E0�Ö7)7_���c���%� ����/az��1�0��������e�t� G�RvF����/�&�2���$�Q�M��(�Qiqc�2;��tD�|��3��nA �IH+�L�4A5§$���T�)̦�5�]"#�R8���^y���K�j �%_.�fg8�ɶ�7��g���AP�}����U���'X30C3��+�Q3�)��*�m+l��&�AZ�ć�{mG��Q0���t(|cI�WzF���=/,��{'������j�C����۸�\�z��\b|���LJ����NL�� 7� �n�Q��y�ps����Z6���;-��-�q�N�^h����7�0ߓ� �J�A�������i�A���a�6�}�rB�h�H:�<}�6������
�a�og�i&���n&s��x@OM U���}��ۃ-G1z;b���=���F�%�^���9�0��ܐ��W�Ǝ���g@�F��ѕ��D��T�#P	,Xv�?2?�u	-ג���[�{�dv��DЎ�Ŀ���k"���]���t���j{������JO�[�m�j��"al���������E4e�R�OY.v����a:���4��^�X_iU�ծ�����)j�f����:[�[2��K�_>���Z� �B�>2����IĶ�nUZ�1L��/,�Z-��!&)�����S�D��[��毾
"�U3%��3t���v9���H��F�ubz�=�)��7��50�Fr�T]�@
7�G�r��"04w�1F�&Dn$�;��:���+.W��*�`6�NԊv`#���Xy��F_
����.�+��ҥ���I����{�U�X1�=�A�UCʽx#*(sG����+B��lo�G���U
Ui�t�x�����h�S���>��(1a�u�����(Π,u��Q5c '��;�:8�V-�L�0����
��ľ1"��Ut��oA�c�&�K���-�4���`o g������rDٜai���-�#I#p��b3s�3{��t3�^��-6xX(��P�Bn�b�c��ɬ��y�s��@��ӫ������%Q�O3/�I/�iLR��bJbE����T?P����������J^y5!���n�%���Շ���`�? *�b����yfc���5��9��a��2Ke�&��o<��i����>'v�4�2F

����m�$mx���H��T�5m}叠�Ax�������5?v�_se�恉�����3ҽ�F�L?7E\m�N"���$��n9�Uk����fu�y��'������o径�K�;R��$�zO���9�c��6w�ؒƕ	<���mI�rn�= 
p�����-�
�u	,ʘ)D����.�� d٧gZ�َ�sf$oN�M��ax��3��X'�ȇ]�jJZ�A�ᝨQoF����7�QG�w���g*����i�T�E ���ς��4�W�2yp��iI2�	��.#�1��,4�7�a����P��"���<���*L���ϞrLw���*�)��Sm�z�K�pS��+��"�lIj�7��i�^#�.Nm�'����͞��Ǧ�Az�s�g*����k!=�:K�9�Y����A��\"�3�5��
p���t�v��b���כ�2Yc_ �.���\���c���ԭ?��f�D9�y���U+��X�M��`8xN�I����|�v&*Y�=F� @� JF\O��-?����G���H�3����/߅"�[�i��H\�0Tn���E'�����EJWC�WzL��C�}Byy��oW��֐R���|d�t=�i�*����=w�_�����L/)0�s�15���ʙV�c��S@�p���l����R����k��sQg��U)�n���#��U�J4h�;E��V���d\�[x�ֈ��a{�}�('+YW+`M$ɓ�;xGi���Xfi�@�@.�>�e׌󛓿{�����_^y3��yv(�����hC<a�3�bf��Z�M�N~�yl��xu_>��r�C��g8���Q.�
�G�yI�B�Gi��� kG���u�c��Yb;)DP\�j �6�|�=�^��~ŀ�ӹ�y�Q�2��ۜ�I�,yH^|&�5���YG�im�5��I�n>`Y�	�מz��@G�::EE�����W'J���(��[NV��Uʃ�3Z9dJ��"xABm�v�F,J�FV����F�q���e�{�r�ؘ\g�h�8Wt��F�Fk�<Z���P��Q,/�(Śk�	uhChԦ�"ӐOh��Z!�c���h��2m� 5����=Ewcb\�At�;�3�^/�����zf�(���Ǣ�����,m�|D��'X���F�G��o��l�����T�wS��v��,����`*�,?��D[�x_�J�f���h�(���n(_��z��S�(�U/o�����d���� �X�wY��; ��5��q���^؃���1{���ƌ�)���>AwFize�'c�<�G���TQ{���T���8NS�� Q��,���Ц�U�w-q�^̉ӧ�g�E`+���D��O9Pفm���;�׼"��?�D9�9d�п5���Ɗ5K���be�h�M20�xG�l0��w�q����j�4��6��I
����L����*˱�C�#6�Ҷ��׃-�������.���`��(��ozC��N�ΗA��*o�d�2[ҥ~�f��H�]s�����hMp5�嫒盧-�$Gi��9lH��-�VU�R�9}�ЄG�I�ZAi��tXoYj��8�cȌT-�h��sĳ� >
wbz����y�K�H�� ��v$�����#e�S���ͭ`hNJoQ��������L<Xf���3d���G�ͣ�!�6;�[�ň��m*@�%��f�?sQ"XS.�P�7�a}�(B�2��0����rR����=K�; �9+6��Ҭ0x���)��u.}�@�_��,>��1�2�Du١� -��f�)䚶�(w�>	|��^�<Y�hw�I>F�οt���f4��\I�Q��W�ߩ-q���+}���l����Z�����]{�UDSq�|E"\�m��_�d��&s�R�1��[Q>�g�;�+18�J�M�_E� (��d=�]q�1ʥh1].-�u��@�Af�h�ͦD��Q*4`�|<�N��m��ᚨdl1���8%]��� B˨�@������I��y�!���Q�;r,�K�Y�u]ݰ�\O�m.lW��ʓcGc�.}��L����h��/�,&P�Y� ���J�C��8n��V�Ɉ�Ҷ��t:e�@����Z�\�k2Y���b�~��UI �+T�_�CP�!;F\�����4�*�ý�+�U�]Kr������DYX+fX���򼦳��lK�5�}�k=r]98؞
\O�kC)�g,;�!������0 ����#�h�2��v���#D��D�b�v��_����p>��n'ɪKA_Hc2x�̃9b���.�1S��u"��M,[xdksh4�W� 'y���.N�U��}^+!s�-mk���%���%��
ѓ���ds�6��� ���Z�*+o���d���`o�����3��|�O�~(��*�~̆����9P�z7�i�$ޑ���%�I�C�\�o�3��(����g|@�}��˛�m>�,�����Թ��f� �L?�r�h��a�M|�z*�B]��r�W
i���!{[�	�"8��e/�FHoI�|ȡ��%U�n+�ŉV����"��9�\fnj�*�.(x�I�NC��5� \jؒ����H�J���j!�������J������Jc^_P�X���m������h�r���ك;as���D�u����gsj���ynpZ�͜�La�5�n�J#X��u���fQ��eTOSd��98�v��.�N�������#�͐�����#,U�?W1@�kAy3 ���T���T&����Wsx.Z� S��.2�,lGV���r��O};���:��Sb(��T�Yx-\� c�����i{�&���Ǆ-%.��	Ɵ��)���<U�M0pT>�K��Nb�����^���O/������y������\n�r�p�Q�߭�g,�c{���21�?+�Rb�k1d�J���*;��+̢Z��ᅵm5ji�B5�&
-(��B�a�t�����/D)ߞ3�a��a?�n����C�j����RgA-u��E�z+�=��A� T*�V�:U�M�u$<���cϹ�P#�����Tz�
���%��y�)U���zƇ��m;�塀�����$a���ן�n�֎�9-���q�Z�R�J�p�2z��e�]�K� w,l�	�*Ⱥ6'M�D	��ޔC�*Ḯ;(�!�1cu`K����m�B�NI-yK[�:vQ���k��JǢ����O���a�&�������,��9�L���V��KQב�7�6�G�5���߾6Ve����/�����]�]�K4bkQ^X�5Q)��1��A�bfa�$*h�MK���B\l�F�ۺ��2D��j����ONb,���Hx��N�?O�2y�m����G�eI6t�������/'���vZm��v]�\b����Ԩ�����KGp~�X܋���i��(
{�a�ګ�_�<���ϙd��i�~2MRط�8�߁h`��|�+Or��mU`�V�ʾϬd!�]�I�L�1�`�z�?������`ƴ{;���B���i"4>Y�Wl�N)�+o_(���|����ro����Υ��7]ű���x
���ɐ5��y�u![����
v%Ht>*݊�37���4Ey��h��L�=A�=Sm�z����O�Ƽ�غ��[d^�~H�R�X��HW�2 e$�n��o�%=�Ҙ�����o�v\�&�*��Z���7�nc��h��'ET	wE%L5�W��lK�HH9�]r����Dn <�U�@���]4U�oS7!j.(TT�O�.�$5Vr��J����	|-R��=E0���%6#g�,��OihD���/$�$�8�T��eg��/�'G���JUwQJIH{��G
�HI����]��#�
���v�������w�;��Ú����J[GZ�r�2����F^�a]�=�-=+q��Dy��I5}�Ly ��َ%����tqC��I�0�0 M�ƕ �RA9�{�Ӯ�i
Uy��J�u�9ׁw��L���҃(is!��������p�#���T�@��bEf�'��:���R�b�0 �8=�.T��k����e�&(wc�B�6�NBk?�΄7�����[n4mk�y��bw�)���,��,�縄�v�q�`HZ��^ꅝ�M�3�Iȱ��{�!��Ѿ~�4�Z��l�a�3��{$l�bsf���{�Kʙ��bK�]5��>����Nh�M��|�_;l�x����u���w�FqL^��A�H��\�a�:]؃3��9�|�n�I@�i��������N,���ÀR�h�/�aG�8_�խ;�a�����6C|���Qڗ��.b�H?��w��|�/�H�"�{����:P����B1[npըH�~nſ��� VL!��i;�4'� bͤ�]��vq{��Pk���wJ��!.�h1C'q-�i-)�C2��ΊӮ���N��6�R��?�S����yc�άq ���f���qT|X�,6t������|��p��şlC���ªE�ϼ�9� _P�I��sU�����/z������rWs� � =�{����������W�[�z&�������2za-�b�$'M>�@���X�)[me��I_�)��q�~V�$�Ȋ*�c*��h���1.r>�,���}��&8���B�4r�������wr�gs�V�%v�'�}0��eҌ������e��6C�}bĞ��^=tɭ�I1�T�?g���)ӟ�EБ��|4�B�����e���^;}���f�+v�Z�#������S�W0�L7e�]���M�$�$(2���;.���ua+H�t����qf��7��_e 1B��+E��ǻ�|J>�=r�!���e�aܨ7	Ԁ�d��V#ܴyBE0~�s���W�e�+�M�J^7)m�R�`��r�W���Ѹ�O�O�/�������;�y'�A���Fi-�T���q�wa2M|Ax��Mmmq����y����;��W�j��eG�#Pd�,P�kdZ����ѷ��.43/,�8{����O�
Ԉ>"�1���@Y�"E|�A�|:���#���(M�4���uw6��n�?�������<�W�̕c��,�{���j5��y�^H"��8��13�uڊ��\��DH=�����B��]3;H�G ?=�R[\�����z���1SdU���u��lr
�\�#�� K�h �xTa����Y㉂I�<(�`�S�H,I7o_����{�x��@�j8-��z�ŋ6���`rT�b���uи���w=���Ɔ	�h��BJS�������	B׬DE�G0��7H�0-?�AAI�_,��;qQ�����/w����beY �r�:���o@=��Ք����`�h�0��Q-H:���@�0k)�G��|���o��9�F-_tS���N�BZ(�T6v lD�h�$o��a�gq�C/B�}z�X�eM)[�'F��k���t[�b�E>� �Ԣ��טE�X�g�\p?�K� �0ς����!Afn����N�|��`�_�-2�x�Eg<���}�0xy�Ի�	�B[���5��1s�A3H��|Tn��A�٦�mG�����	���OM���.�� L��|k� ���j!u�^Ra���X�L3��y�4hV6�YPc.�M;��q��^�uv+���ҩ*t��9�������I����O�]�mn�[�1:����h��m7�Ld��̟ͬ)�%"c,�j��m����0��{���^�V� ѧ^�5�����[�vI�BK���<G�QD����j��큖N��5,0ܶ;�c>�A�x���h�t\Rh��0�8���EcX\��G*�|�-���v0+�{,��%]v���s���Ma�f�~M�/�+O �'6�P��a3>���H8�����r������e�����R�%�<;+�q�%����&}T����5	ԗ�s1T2ZĘ�R�I���u��7$��܅�]$��6�V��Nvb<���%F#wlA܈����!z�u�\��`�J��!3�9I(E?���/cq�c$�	Ѐ�t��w=�x�ڰCv���D:����f`�m�7���(�*
+f	+��e�ߥ�1`Ę���m�::��r?��(���S�����4=��SD���� j[�&�_���M��xY�(���c�ӕO%s�ő�tt^(�l
��]��
�u$zW� P�B͔;_<b������l���O��2��s�g��MF2��j���O�4	e� "[p��W_�K)��*y,RۅR�����fi	����sd�F61��!���`h�u�����doX�u���K��r��Ka�G0���.1��#�8I��-�����fUy��J!� ���0J�,�����~�g�����(6�Ľ�@Y&f03@ [6�� H����k�-�G�#l�	�:
�Q�MN�$xp츚��p@��j�Wԝ�Z[I���>�/e q{u�������}/��zJ��@�9�z2
�8��1*,3�eqZ��� B�� ���C��x)��^��w�?*p��`y����	c	;���wї�^�qF0P�<9��0�.�M�ASvg�{�ʙ���p���`��Z��62Q��	RXm8qC�,
-��h9C����Z�- h�ؓ>qH:�.H���1����8�:�\���!���%��c��wg�Xq�	`T@s��lOA%�?u�R[�w�DK�v!��M�e�f2+5��8Рro��AӀ��tTaH}��v�p�����,�P{�=�G���F(%b�����F6D��
r������r�q��>��2m}��U=����z���p5���ssC`l�p�e����nE�c'�K�>�d9��,��z?�Uϰ����:�҄���q.5���Q�T�Gj/�XC�Mc��$����Io;�R��*vAeߴ���Zy���rAz�����J/��rl�������9�c�
�%�(�Z�:(���m�$��W�V�so�`��Ct)z��3���慂��/��{�0dxk�a���sfZ����l���Ů,��{�'���>����+:��_zl&7��f��<�{�p`%.����x��������e�zl�c����b̎-'��<�{��\��.��߉�����
�_SR���Ρ+y��nY�$��_ٲڕ�2�\�G��B���fC�rgm�v���C7���{-aݮ�(�N�s)�;�I��'t�AN�?qOB���&��1`q�S��ˬa�7�M2O�'hv� ��s�E�^�R��A� Ln��Sm:B�Y�`���Rn�ч��%u+;����\�s�,i�(�6Y�CGUz�n��S$����xP�_��Y�*��:0�^oٱ���\�C%؈w4��q���m"���?i/H[P���P���I�]\&�)�~y2N]w����FJ���C�T��0�V�(�l�@��1�a,NL�@��a��͋��V�z�f��
�[��|UOܻĤ;�� �C@�� �쵘c�+]�kA���:a��77�ܶF��T�Ϭ{�V6>�raZ�Vty��(�9�C�RS
0rSC_�u�̄ !O�[����?¬�&��5�Pǘ��ֺݛݼQk4�w�����t����0��{/ �; �1!(��ܗ�^Y����a�vǅ��ZyoÇ�����נ9W�k�xjz�U3ǖe3dDk-w&��<�B�-:�O�{O����w�{x��!ű)HqDuo8|r�b�5oTLq?�2adnB�Z�����3�~�"�z����ࡆ< �����Kx$`.� �UۆCo>R��1�~]Bz��Zƞx�Aq���]��A��{X�̡}�e�ȵ��ߓ���rq#g�6Y�GP)��� <s�2J���cR�+Jxʳ�)�hk��٫�(!�ԧ׳�ʡ6����&̗�"�ӻ ��P��>�0�������J-��D! �,�*��(}�ċ�S��{�׻0FGۍ�-f@�E��U}(�������{�C:<8uO�q.�G�T��I��D�֒3K���KP����,]�#�X�� ��س�8�����p�,��UB��B��Q�@��#G��L�υ�O
���	��C���������V�f8z�Fފ�ؕ�����KC�$+Q�$��Hz��p�o \�L�b#
baZd`���6��.QKSTԄ��tg�IFA�ߓ駛դ_�����X�i��FAy��X/_�Z��rn��2�aOh�iȠ�!
D ��U��_��>������Go=Qp���f���z�����=)m�cd�s0��-C߼A�m�""��ӷox��ڬ&U�R���_,�4���'�U�{�}�Y��"I��[8��*�"�6g�t�87���Jgv$�X�-��ڍ���l�����a&�Sa�'��3�B&�r+�&]i��8K[ӞΥT~�j�mŷM �o.ˀn��3�3V{��T�0�];F&#VW�^t3��r&�U��G!��}��#��V-m����r@�R1�2}h�0q��{���6��0b�T�R&����@�ZO-1m>�o���"�is��ૅ���]+�j�'$H��p<B=��A3�Wۣ�,�NxD'\6C�����>"
�~G�]֞޽+0��FG_je��w�Ľ"x��c���k��$H�r���<�9N�}�jL�5�I0��߄���u��c��6�簶�	��{Yۯ���\5ϜK��*�d��,_{�׈�����ߑ���d�8�m��acX(�rB;9{$,�J�bb����۶�.=:
e�P�5��z	�(���Q��H[��a6#.�6����f+B{1���?�m��,ꂒ+m��U�Ћ��o����0C� Bs>>�������$EHf^�N�#��sv[�
BXծ�h<9�t+5 ��c�g3*.�I����Rc�x����|V��`��U��o����1u�	����C5�Q~�oz�a��2��e턈c��l`�<O�#T�lɍ���J��M���vp��^��߲��R<�q*�7ϳ�L��	O�Rg�f+��3��[{I,o�D�Sܑ��LB�B�� �-T����X��¬�ۦ��|}��l� #�z��}����q�+������(D�6�S~Љ����<M�tU�6:<�#�l&��3<�߲�������	|�gm���K�~�T��;B8XS1���w����>� �2"T�����y(�I!�EJ�U]�!����m`k9���rc���Sj�v�����HІן�_Ѱ^��9Y�&�:��U ���E�S#^��Fq���rqIkl?�p�P�ۇN]�U�ςF;�\��]��+33����:�� ��͟Ci�g&�&�LQ��r���&��_m��ZXW�����<��)��u�OqwW��?t+�70�P�0?�N�j��E��[���3�_Υ�,ɗ�TZ�x����/<y��@��5��w��~�M�֫_���f�9���QF��Ć:BG(^�5G�:��"!����bq�l8�Cp='C	U�(-HL�	V�ܠ�1����Aj>�F�ɕ�a�����sj��X����h̜xjx+_M���V^�'|��Z|��C:������(uء��l-�s�k��E��O6c3��`����C_q��?�C���J_١8B0�2�m(�s������eag�w�E��b���u����(.�(n�Z�|����h��DO4�d��͑֐���#yN�IM2�ѓ^��}��X'������X�}]<PY��Áԓ?��#���w�]���Ff�s;������A��鲈w��)�����(�����5:���t큮�7%+� �Q6ni�_�}���īOT��)4*�o?�I��H7��}��V������{��)M�`�E�Mx���yBB�a�� %�Y�N�P���� �߇�s�A�o��g��_�V�&v�A���K����>�j.k�����_u\J��~B���J�6�X�!�����>��IjY�lF�T�n�9;��_�RG=�@���o���:�
��Vd�=oxm���65�/�[���HjR��k�?���w�+A)j��YGD�1�6o���=@Y��e�D��Jhy���C�־q�}��)C�ѸW�� ;s�p�-�t�txn�]yU�ߋ�x���1�b+I�,��zU��Gv|^�P�m�_>��)�X���k�2���ap���!�1��Z�uŃ�w���#T���OIy�]����5����_����P1l��J&�Y<�[�����2~<�<�vϚ��a� p��j��2"�ߍg��B6�&����!$�.�C�O��C�|C�L�@��w�y�+�}��ý�����qR�Q^5X�P���J\�Qn��trM��ؐ��8;Q�����K)�a�����CA�^�g9��x���q3���M:&~�髒Gpd�W{3�����s�o�t�Q��#<}X�D������4j�\�р19
VHn��K�PvT����b�~���nTT�%U�7>�n��&#�%����6�U:*e}&.���B�9���yA<D;(k9y��N�/�	�ȓ8c_N�2l��[�gНr��j�a��� 6�N��B�
��ɴK/�D쎲�<�[o���O;Q������Ԓ�o>=��ǖ�`m�V�zn'�.Y$|��[ǧg��ϲ9 X��o�/���r5F�A`�t�@
���w�	QW�q�����1�@���M��<���$����M��%��|��M1 ����]���)��~Pi��l0m�n�l�@�Jd�w/�Y2%h�kR���#MCh%�v
-WN�t׵�vd��R=��2wb�N%��m"!�b{Q�ߚj��ӵ��{���9�]�$nE�$������e�q�B$t�����vH�
Y�m}g_���>�dH���3Tu�Ѡ-gk���u|���0\MM���˭W���H��� �����f*��[h%ɰd���#���#�T�q_�$���$W�H�m�>���!H����O_�Ԍ��J%ϸ��C������e��Ɇ��G�Õb��䵚i������ռQ�^c�vr�|���I���9�����3�0%Y�A�X�{�'L�g0�ܟR���[x����g贯���eniB�L��X)��Sե�Ikǽ�-�$ǝ䨸���,�tLS,��@/��}�"��>��T\M�[�eE�j&��m���|���M֙W���gtt)�%i��E�l���������*�8B����$;g";��;�N��d�wywN�,���2���|���{'�K�a��&~�5��dğ�����R�ÖC=�׆�X
���"+~���hu'W��oQ^�$UV��yỏۘc���,�cycKI�ʂ���Xia�2��J�׈�s/NV@��s�ӯ�}U���	�4,嫁�+(9�z���[J�vp0N�Ы^]�A�OI�$T�<��8L��`��S�M�D�o���e,��ֻ*�X � a�ZY��������1�:uk
���E����$�m���OJ�9]n,'�%�����U��Ɵ�
$�Do�@�JX{��)g�7�� ����{�K���k�5�\������Ό�DC������Cچ���l����m��	�o�M;!���0HWu�vZ�_��4vZU�אT�D�gWL��Jk����NL�o#5-*��X@*Gz|�Eu�������	W���ϕ<٬�-ݹ2���<ǚ{2�<���_�;]lʟ=�z����y��ൌ�k��ڌI .P��
�\.�14���ݻ�����+�s!���H0̝|ʟ�Q��r�*s~���m6�<l!0�ŝ�ko�\m�>�	��⵵R�ϖ~
��<P����n��eS�Z���Ojcl����h����9�h�K)�Q?Q�J���5Q�mD5����U��H�D(ϭ�ؠ��ϲ��uQ��{F�vr�#�h�8�<�SJ�@o���ٟ��8F�|'0�rEưz�Թ�H��Q���m���[]���yP��/�����\�%W]�^��E�*h?��@��cE-�h��xtxO3i�(ޠ���1H��/5�б!6N�
��(�>__�O���{\�.�uՌ�����yk�	a����Y���H���הL�Ec�d ����S�za��@=W�!�BI �S�>82D��X�K�	9[*r�ˎ{����~e'��e�gv�0���Z��1��d�F(�$�+D@�(L�⒦�k��Z��[��G�� ���(�Ů,y��m���\�^���)�2��6ߊ�]�0���]ۢ������b	A�-ְ.����S��q�N���,��%������?	��z���(�K­������#=ڜM���48�?�Z���V�/Ejd
����E�L@�w� s����U��3Pб��Q�z�����
b�(@Ez`׀�
!IV%l� $e�2M���E����
��F��{��T�jH��j�7.,������G��SIJ��÷J�'Xo0�]��#xK*�W�K�##P�f-�5��M\_U�(�iW�Lڢ[�]c�%�T�T�__�nJ����T�H��_�4���������_.�?��s[%}/@��8��V��е��G;���Cp2g��W�(b5��S4�gj�o�$��ߧ]>�8Q��O_v�~�����X-�\Hy�|lf��.��6mQ��iz�O�'�~�D�$�����_��Ԧ4�3ui�#��u	mO��N`�����b�&��؈\1h�-W�����ak�G~y�2�ȤФ(�ŚD��&5�p�Q��7���`��s4�cM�>�ěD�� �̯��jd��;?#�	�8_����$�'���������hgzRNLˢA�T�˖�zsax�bA�
�YA<�01�]��ۦ��1 �A��y>�>x&�&6�"��[N��d@�߽�"P�t�kZ�[m����[���r+yxPy��:Wn��IY��I�́`<�f5�����fA�n����w�.mb�\ƖrerC�C���~"�i ���`Ka���o�G��_��/��F���Ȫz����j�2F�y��.�����n5���8��'�lc�^O�0�đ�����\a�w�-M����敥��!Ϟ�P<��8��%~'��
���n)ު��Π�b	���,�Rl��	�����˧ph��ӌ\8����5������P�S�� �z�&M7���u�F���]��RP�U0�n��jH���D(h��r����J'gj��SeW1e�"�h��J�u����Nc�u�s��琓�y�+ ��q�Z�(���ˠ��c���*���8��)�qo�
p��X��Z�sȮ<'lHT��)+$�M�����?9:g�D��"��h���Bv�:����N.|Pꛖ�:G�	��I�\���C��>���0��eT[�R�hyrٖW�+4�b8�+M[(z��RC��?�\JV�N���� +Z���������%��
T��l��U��rP{:����zI
4!���~��W���9���(���H)s_��ږC�o�C�$E4]
(������t�SD<�rӃ��ޮ��-h�7v���v���i��X�=9΋��� 	�F�b��'['�ȏh�q؅7ͅ���([+p� ſ� ��:x���*i޹6�s%�i�N�'0׵ʓ�=���`w+-z�̑1րp�J��)�v<�N��.�\��|�j}l�B�5n:�ET'�K~�+�N	ŞIӞR��{��J�r�P}�^c�S3�I�S�����u�-����CM%3)����Ͻ.l��zji�n?Dy�,}�B9kV|�AqFoP�UytU���]������:diVtDvc��00P��sE��6D�����ٞ�(���F�i�݈�ƿo-#��f�$�ն�ʹ|���T��MT1瀚TZ:��95�9m��6�'-� |i���q��$�P�HI������F�<7	�%m����Ӛ���c�.��'N+9L�7G��")<����2|����de���V�����������b��g����0� 	i���91l�ղ�����3όQ��=�m�f?����TI��l(Tl��}ϠYj��XS������q��y2~�u}�T}�$��U��'��e�_�	$����;!��p��w�v[�؇�z����l�H��Q��C[���ϐ�� ��2���*��{�]5H�D�P'��B*�M,UZ\���5	Se��?n�5�o�
C����rL�Wk���gh��ym��3��c_���f:�H
`�t=����N��:M��&�U��)[�����}�ݪ��c����Bw�$��*��Znq��,|g�������"w���B�� ;�@Yp����g3]R+� i�_%�f��ܠ��H?N邺�o���*n�<}9�oo�����*2��T�k�"2���UB"F���Qo�W���������Q�|Ǘ=�Y��9��|a�9�C�֝��/�l�B��K.��M�<�����9�,*@�7-���ET i	L�#�D&��"��ȁh6�=Q�7ŀ�gY�i��,��:V��VwA�Ws�{�ΙQNCYF�h�0!�r�P��-��8������q$�"�9ѕ?{��F��<����G'�Ū�u�4+e�+~m����2�@�Ѡ��^��Я͝��&��%��HQ�R�*Y��7�e� ���W\�]/�гi	�QH��c�
�ߝ�t��F���Ȓ@y�S�?��^N,g��"��I��7�����~_�m���~c(���v��^׾ߵ�8R��@Ó�q���V��Pֻ��~{����xۃ�V�A(z�d��[��,���}�e���Y�j�_�����&��^��:^ �[��a�J�W	���$�]L�a0$��EJ}���U-��m�z�<�~�1%]�EH���\[�䐵��>��Wg�l�P�Ut��c�2�|e\h�=C�]���z����3 F>V�|~�jm�`0U����t�,�v�ȝӁ�g[v����}%���i�jbn)�?�� �?��T.��^Y~������_N&��+(!i�������jsLC��zRTSw�U�� �$�2:sۿ��o�&����`�^+e$k5��'�Fzw.��Z���X���T-I�#�D՟�D�!���|)=�PJJ�Nt�p��<^F�9���|�jУ��*,��u���H�Y������I�@�1G �}8>���t�����$$3�Z:���>V*aؓ���I5�����Wi�<Ԏ?��L�q��M4��ztD�����H.��s��3��s�4]  �D�T���3}�xX��im���0���!.�Q0&�kݤp"EV�b�Ԅd��p�f�\Q������� a2�[���>Qc�QG0���1 5�=�e�ւ���e�3�Fɧ���MU��L-����:Vo	x�K�z�^�~�."JdLc*B����]���˽��U��O6�l�}�`�,��x[K�ȇZu�ϦU�
��f�b��>fˈ2~\�4Tg*�ؑ.N9U�0�U��
noj�ͨRB�B�U|�褤jT�λ��%m+�ם���=W�bWK�%'�煍6�#�Z��?v��pvn�D����K*nS�.g����u��#}m�%<�ϞLI�����P����&1a)6jOt�!H�q��j��Z+����c{����L@|d��{���@C=��mQ�P���\t�{�<�#�q��k+_��L@�U��O�7F8DL��AF�b�����5"���C4w�����A�V�C���(3�	dUXߎ�K>����e"�}�x�uk��iG;<�W8^�ϕ�ɯ�H��&��8�o����qIucM�� <�\���'�V��������+�Z&�Mz/BzI:M.�3�tD�q/&'>%�<�������l��*�O�u����܈c�|1�4��j��A�Bش�>�e�^���KL��|R�)^�#F�����&�UV@<�HT�P;���ѿ&�cW�l^�d� �<,L��6��'��eќՃ�Ҥ�"���:D��#�Q?RI˖�H��y�nK���V���|�������F����j Pr<��9e���˫F\�e�Q@f;���zL�Z4�z	[���m=yj9����؏u�"���q��T��5\ ����b�P�nT�PG���x�>U#����}�F���j|���6���>z���uri�����ִ�]�c�͢�k��*!�h��J`%A��߲r:\a� ��������LO[{��	�u�&5I܉�BC�`z��aZ���1��	\�;.��1�R�|�Ϸ��~��(�#��T�d�"!�㔋���*����쀞9���z�F�?!Y۰Y-��$b��1m��U�����N� ��NǮ�V�e�C��9?J(u���P<(�o��:�{,6��2f�켢ZH�]����l�ɘ-���¡�]����.8)Cɏ]���<ЎF�O,ܔ)�B�A5�=⁄Cy��U�vW �9l��%Z_(E55`��3�D��U��63���@���h/��t�Pm^����nߊ�nA��xr��^�ts��F�uȿ��`u���w@�i���\��d ���u����������N�؍}�[xM�;��$���k�O��9��?У�3=	�����A���$hP��S#D�p�"��ĵL{4�rzqѫ�BMօZ��*
�^r���lx������}tPA�4�E�"�
"Y]���|ߒ樰F&�/ـ\��g7�ʷ��J���b:!�O��Mv;$�+K�;r� 6>���V	��f"�b3p��|�s1n��Y˲�J5uϨK�O� �7.�P�����տ\bqӱf��/��v���@��+�㣱a�a��,�Q���WX��q�3���Z+���e4�B����1�!i�l��숖M"�%8V�*p�@ԤjB�� `�O:D����Y�Ҕ 1��n�
~��N�\PW+��;>���ͳJ[D��y}���Z�qY��km���Kd7��/�T����b�Q�i�}d���\���.*�+�%7tC�싷��E��Cl�J�:C1���G���6��'��n����MM�ȧ�e�І4pSC�zf�����X��X�B�(8;���(o��±|4-=I�P�p���V�{)��MO3��#GAkG%� �(|�~�k��z����P����-���VQkP��z����H��$��8m���J�;Ag�_�ul
*��)��j�l�P ���p_N`���UOkJ��:�Z�`?����R��3*F�Z���9�Z䚁M��ݱa�;zb�~���N� �Ү�!��d�IX��^E����<�*�* �N�% �5$49�C/�� ��u��d`@�Ld�u�#��� n���Ō��06�4Yp��S_��)~���>�4��P�Uf,x�"��C�c�g���Vy�G]�|Ӏ�H�p�#�oSVy�<��ל�@ł�%!� �-R�2I��P�q���.Ɋ��pFG=ø<q.?�x�^0���(]��Kp�X����7��?�ַnM���k��n_�J��w~5Ӯz�f�=T5�w��!�a�4̓3�5ѽ�T������#9����L�M���f�x'�[@5�X�'�o�0ܳ���ٕ�R��z��FYRLq��q�=�,���Jh�Yw���M�%Iº�\�`[zB���Y�ԧҳ���F!�˭���cZ3$�$>JAC����Y�*ifF��푯�F{���<[���K ����E�~���.}�ׯk���
0�X���<k�[��W�Nve�jД��A��ؿ���t�����/nsGˀnH~�S���v����Bsۮ�����,�$�-���;�c�����V;Ί%R����ޕ�I���r��O����S�Uԯ�n)A�~M������b�S~;��v���a1�S��ةa��bQN\��'�>��tO���B��1�}�P;5vd�t�lJi��u���L�ɠ$"1���4����4�͘5�=��x^p�����-,��AZI�q���w��ݖ��Vs-5���s�$6a��ċ��O�!/�'�[U�S0 ��Ƴ��e ��-y��;���Zc;O<���Xx1[Vl�'�q]��cw���K?rdB���U�Q��	=bG�6]n8�ܨ���ҡ���ў��Bk�='��RͩO�r�]�.�t�j��~|}��}¿^���+����,D��Z�{�X
�6.��)q�T^�E��[�}����_U�?PS܊^�R�̀T��2�:���w@֥��J�w��m<K
��2�"� ��;��^#��FA�1]�4�*03�� 1P*��?�gb6Fgp.��,:�6�n��~����sݢ1��[�x��+��%}P^<&$��d�<�����W�ґ�괤6:�����u0y; c�G�͘4���	)�����a��@��MnQ6�6kɆ�b�s������J�\_e�_�f#h�Ig0p��ǖ�cC6[]]Y"��L�,�~i2��D��uA����[�sӊ쬯�'���$��Q-H�]�Eq%r�����̵�^�j ��י6��з�Iq�X��J�=��?��0X�j8���J�Wt�A�?:\�[��|��1Yȁ���O��P"*-g��{3$��ߗ�~36�p��!w��)��y v�)�u�Z�'�N3��1��=dA��l{L�J}�`svd��EQ@��YDD`�½X)ŁH_�� o��  �%���h+��;�V3X����Fp��/0+atH-1u~����ߢ����iV
+����vv��*&�3�4ڹ��ɍ��D
��y�R��+Oۛ8��0m쫚�����1H`w.�QYR���2>��VO�G߸/��Q�w�_ض�E��@�6�����%���"u;��/*a��-�_.�����7]a���%��M�����`7�Ȱ\��5�a���:p�9.GsRt����m�P�b��TP�P���:�ea�K��iE��U�c�[KQF�,N�4�ľ#̆j�G��[�$ޕ�܈3W�,Q�>F�g�vO��F�����޿��K�T�v�E2j�+���9�񉩺sZ�S;hnSMN4Ƃ�\��[�r(�IW{��|�l G��v��O�.n���
M�s��s`���8d,��,���&��v�Q��o(a�J�3FY�!wre��A��?뙫�goۮ�ݮx���������fMm��Ln�R��)�z�!�R1
�c��������C�)�Z$~�R5_?�d�h�_�#�v�����l��(�&�b�iPhˮ"�k���m�H��+�Y�`�S�z(��#�T�=b@���~��D:ݸfCE�q��X�6�BՅ�V湰
r��VHԶݗi��I��z5gB4���, ������n�T��PQ�����,%�TG7N��9A�}B�N� S[�b(�ޏם�]�#�Q��;��0�οlɾ�b�Y���2#��[�x6ܣ��,�m�T���χm�T�0L3l/	�-���o��>[� �2��UǷ[��6���pى���_B����T(<*9��YV�kȓ������r]7�oޙ�H� 4��Vlg?x}���m�f�ܜ��W�������/û9���M=����n�o�	���O�{��=�݀����Z��_}����2'*�pJ%��� {uZ�D ��ݗ��2�����rY5ai�NV��)+��4L/�é��Ovj��e�$_����v��{��~�x���Z
�J.Ǎ�\��#�?I.Z��hڦ�B�E�b' ��Qǧ�s�qf4���LHc�8P��VX��,V��5\���5�8j���vq��q��Kn�oUzo���#�5l�.�L$Xp�l_	��fТ�Pm���N�N5�`!nj;�ȃ�0Z`2���l�.��ʤ2Ǵ8��o�'})�a(����_�2����� ��F� ��z�y5{��`X�%i�(91�]�Ջ:��-��I5X7F��BJ��&X�`�{}��>4GыX|X� ��X�z5?��݀�Zrkd�U^��4�9"�<����Z���˚�����u�9w� ��w��B�w��H�����>&���E�|&�ߜz&f�����1��x��W�
�O��f=���\����&-F�ڥ�[-@����8,�: þ�Q�f�݇$]�a�{�ghtƾdb�J�	��"D�Zݕ�y�e�E�.ax�K�uW��ݨ(���w+��	Xތ��uU�P>U��${��r�$�l��Ιa��x�S���+�e��NHI�@�O��iI/��w�wfҨ?D��M�i�m<�Hy.P!\�U����9m�x�.��#8}�� �D|�:T:oT�t�����ޡ�z����d�ޔ�W����SL�z��-R�띟���e|��^$8�P���z�����G'M����T �|Ԑ�m���9� ��P	�B,;��z�6��Hӗ!���tC�c+g���{~ɡ����o�
������H@6�lV�G5�4ġ�+z/a��(Dɍ�n�����6>�R�j���ݬڎ�C��躚�N�{'@�$0� [��#K����tǩ�ׅ���~�1����%�d���qõ��`��W1������)F��3����I	�EIy{���}�2b�@��&B�"��j��u=��ضL����дL:��aF�Q[���l�5���>�BEg �odgBV�ɤ��`�AF�@�_o���M���U.\��J�-@<x�>��w�a]�+��fH�V�l_;���Ӕ;��p9�d���	��[����O�������fAa�*����`\��|��'�{���}=��+���=�C �O~��Wy�I�k�o�>���Pk����!�5�x�+���Y���Is��B��D�g�?�z����=|��J��z��ۦ�u�������I̾�P���V��-�V.{��"�*��M�B���һ�F�8���h��ۙh6����Ȣg�̘��Ļ�w=t-�8�t:�$l���3���y��X�e����v�^K���Q��L��3ߧ�-Y�v�㨢�nN6NN�۹�����#v�IM�O"<����X�,H�6܊�QJW�&ܠ�̑C��	Y��`3�
�@�t���L԰?��{.+�*�-#���ɤhJ[�T�Y �nՖ��E"�;����Ow�U�C_6��G���c�q�m]�l|[�JH�VIY#x��W��>�5;�0<�>���&�'A�m�M�ԉ�d2���|W���q7>f2Tު2>�����F�!Ų��h ����sP�w�����Uʘ�S�-�5:��a5z���d$�T���~u�:@;o�x��W����j�]�[5s���@a�v�bh��q;o�V�	7F�Jd}̒W�'#�%�mP��Ɲ�x�l��N��3S��NO�>YX�.?qŋ`��F^&<v��w�Aو�5_���/w{�Wrh�Ǽ����f�>;>�Z�����p\�4��<�?�B���^O$@B�"�6x���9l{acB9{�?LSmjA�ܹ]ڠ�]̽t!>�)�v1�w�,1᷶!����G~zn�q�*���Q�<c��I�8i�M:+p=����'���L�T/k�O�8>�wi��Z�*��r���h&�GKU�����L�s���"��[�O���͏��,^1A���L��t����o�Ȇh�[X�tj�	��*M��~�STF{r��t]Ȳ��UW��� =�M��n�)l��>xE��l �\�I�-Ƀ�H�nfs��I;�BB+ɥ9�k콟H�H{'l�X�kw�*0�ex�4��s�� xX0��s��͜�1��Hʯ����1��"����a9x�Nf6�EY�̉Ǎ���If�RZwf��F�o0�cV `a~q5wPW3S��ou��5zG?v�ы�6Zj�����tf��e|���\co�me��w}S4FG�ʆK&�	A6�i��T G�q�nL�,��}���
z#�J��'?Tl�<�J�f��4%��sY$�����
�_��S��J'�R���94'7ё��H
	���C�v#u�����U��&y���|����ҟ}h
h��-��\��c1���v��!��6��y�&�@H`�a�qx��v�fAX���N�Df&�i�g.],�!���>I4���,NP�* �0�H>3��˃���Oo_�R���mV�����Ag�m���Dgo올�b��L�Rth�ؚ�v��4kK����1��t��S��f3���d�~Ӄ��t)�hɥ2Ncwx�Mo�oOZp:�}�iz=B�Pu���G!��P�M0T�.��Fp��O�h)*C�097��plt��ӲK;ݘp�s��8�F(O�׉���;E������f=7�xd�A�߉g��H\ͧ�~��N���0a6n8����^����-F6v����+��c,8:Fǃ� }Җ�V�-�U�� LL���mec�^(6Ly3U����6ُ_,���*�H��������P7�� �3tB��B0���I������zU�.E�m�<��q�_.�"5r����Ay{|h�e�7�q` 8!C��&���s2S�������KČ5�̫�H��4����=Lmz1��F@G�(����lu,�)k�O��up�l71U�~�ź����$�L���|���x/�p��m�o2}n�"��="�`{a�.Kz�����t>�--#�����T�	�?�a#�l�{j��s�Z�ai�iQQ���%L�.n�s�K�?�S����h�K�=��{/��V��s1Į������R�/����I/�	���˘Ą$�����C���`b�z��F�*/HcHe��.&(�ڹ����v�?l�:��<�3a�PMZ�`L����d��~��\3��9�9q�/s�>�
�ڌp���R��Z �����ks9Q)�  an���q
[ݮ�^:_aH���J�����;�$!˘�<��&�=ϹkU�Xh+�����9s���
Q ���{4�M� �8J�����4 TQ�}_��-*�"��ǌ��p=����� +��� pv�%�����ОA�dd�a p�N��L	����"�3�q��#���g�����ʎ�s�՜}#�(�������E�RL'�2����U �V��&ONfuwM=����J��V"u������l���G����e�H�=sH�6�7�B�3P^�2�9� �>�ͮND���^��E�0��bzi�	� �+�fL�E��ؖ�GM���MU���^
��C7S·��\U�`cl�[n��S��4]d�?���n�N^��րX�iG����~K�3�gF*�
0L������v����T�f�����T|��F��lE�cy��ɪ5i�Oe���Xn`�����=�������^�%D��:wUa�H��Q���$�E�U0d���+�G��"w:�c�$-��v�-��t��|*t�c�̮X4�"��H ���M�����h[�|9v�g:�WŲ�.ሑxB2T	�.E�I�V����O���x�"вuo�ޣ[�`����9���?���P���2�����2������W���Lj��˧���'z��صw����?n��Nd���n7�(]a�
���`A�4�g'�kK��I&[���
�E6��^�4Ote���һ��K�}���f�_�9��A��h�5�WcJ�]Y�)U�.$�m��0�1����sJ[�>yn@���ݽP�2/.t)��[G�^�/\{�c6u��/g�\�!��BEvl���Z`<�
x�t���L�`p~�@��!Bl/�?'_�TZC���e7\ ��!B��J�M��a��F�Y�4g�S0T'I2��M�D�A��v�A��ט#.@�C[�H��@A��Y��B�x�~F��)5�N\�
����p~�İ�Yo��"Ә�;������D�
Xk��jsνT�]z�D�(� ?lPd���F�62�8�s��#l{�I��kQ��b�p���+PѢ��-��:71�wCf���a!vb����}��J`5�V����l��=�ICI�D�e��;{�7O/h~�J�i�!`($��GC+c��}f��]/>�K�k�ɇ����k�P�g�m^zyF��H�T�����(��{�-0��+XGj7[ޢ��<�i�g�!���{�����$F�]���W�%��v�:+[�H%�n	۵�Ù�s#��9�Na����h��ӂ �6D���Giz�_�[�Ö�2>�j^�c�YJO�4������$�{.���f�M����v*�E��υf����t�(�ed
^�3�`��� ��ZS�c�����B��_�E$S�=}|zy�A~UD@�OLѷ�i���+qg�X5�n�V�H_���Jb���~�zO/j���=���8aC�HRYj��8�(�3��M�Ҵ�h:�Aq\h7��ǂpV�Jk�_;�J�}�2뻵v��9V�v��/�J�=�����p�7�5+I��}�h�Ě_���J�"q�G	�&1�O�WY��܈�BƵ�����N���cQ���Q%��81��N��Ѿ.�.�It��~�q�|kԞ�1�*a�׏$��sg~Rnh�Z�M`�i��A"��@�1Z��w̓S?��Г~�ܿ�a*w�A?pSz��i�+�*�|��e��4�u������x���P�t�{s�9Z/������/��)���Dt�b��(F� �H0lϜ~��]͊�-}.�D�A�=ղ����<f���N͔�ъ����"����+���e�R�ȍ��:��B�k�x9���-�(�&rpce	s���|[�����O�<۶�8���@)��)~�+'���ǀ˓O�FЃ��¦Q�|e���L]�nF�$7v���"��8��E��!~�y΁����H���l���x�������'z�������U8����,x��)q+n��8�q�F���;���\�sM[�S��IQ>��G� �,E�1�����u����K-�q��=��1�Z�Kp����Nּw�[�����ц`p��Ȍ �A�; P]M���ݫ�>V�Y���}��^�?	c��J� ?	��D�3G񠤴���S�o�-|����_�	�P�tg��c�����+%U��g{}|'˾`yE2z+!]&`�f{LQk*�T��7yj��"�e+2o��K�U@�0�0���0V6A�S��B̑���N��fΦk��={}E�ϳ۪�z�oJ� .�[$�u�8���B�5��E��Ç�vhc)�{�� ���.�oe���ě��N�܊��d�2�nXffj ��c��B��S��'��\�#ߺ�+i
Q���Ƨ�&��څ)�?��ᐉ搵�z���/���4��8I1�����*�#L^���7ٲTԞM~25æ�xP�� �$d��I(a>�E-۰J�s�D*<�Ӥ�^�?QƋQYމ���L^C��O�ރ|���LlG�ͤjf�Z��]�}X�sR��F����k^�%*_���Z��Z����Ж�H5U*FW���j�K}?����+����ո�b�e-��(��;��1@�ۤ1
���'7|{`a[�ZW�Ø�]z�	�H���<O\��ɻU�*�t`B�pz��K�ҍ�^��L�aK$y�>CV�Ӿ,�C|䋿S��h��T�S*������9�$��I�<�N� �1��a�� �|���K�Z�����":�V.r)�rW�·��)��;*�
h^�K�g3<>��'I̟���*~%�ȝ�1�m@��-��;h�� �,.>cEcx�;�����&>̏2�j��|���߅v$}�&T[��8��Hpq���A�W�?x�x�0^����d�=��d̒J�25_[	N����z�s�,:�������y�$k��*S���G�C��M�H2�|���1]����m-��'As9Z�}Զo8����������Š�5
J��?����M[a/!��8 9�c��r�n�hC��No�[T�gĴ߁�jwzT�v��n�C^dT�M��]���n1Es��i�r��NT����Sq��� �ѫ;x��R�F�v$���.wߜ�J翼��Y^C�n)���<�|K` ʂ=Ұ#���Nc �g́$^�����!�M\gU�~��Ι�d&���ݱ�	�#�]3�p�jSU�f�љ��݀�E�(������}ޥcF^'
� ��g���Β�K����Q���`�䁶�3%��=Ǭ8�U�	,V*ShC�}��r9�) dE�}סߡ�!��U���4�%u'(��8����y�H�nܢ������)�+Ŭ�F��J���$�Z��NQ�?SqL���gV2ۻ�ߚ�?���3�s���ڠ4����ͣ���M1��G��8G�|:­<=XLUh�DS�Qi�5�	�a�c�V��	��D��L-��c�����Ћr��\H|�z�=�8Sb92cL���#yPIٖR�Ow�!�S]ڹG����L7b����i���v%NmkXF;-�"-����E��Gӳ#���N$<
���^�����O<�yh9H �g+KU<=�!�u����	��>We-d Դ
Q���2��?��j���}�ÎJ
DT09#��O$f�Tp�M��>^Qᙡ_`V�/�|��)�����4$��ǭ�&E_?Z�.U��LN��m�{���
���0kt�)&4J�� �A�=m�&��C��Z��  �K���=�:����heOw���(E\:�����n	�í5���ܾ�������v�8�N����R��F�t�_A��d�
2�2�t�x" |�x!��Xf���+닡E�/d3���܇/��gs��P$WҐ
v"����b�r�&�| k�M�(�l*���6g�E-�*�E�Wk�r��5T�ۼ��U�O?i��SU�K�,
�y���~=�0�i�T�oDk �O�<4�Ç��g��O��b�K	dH���{;͑6ozȩ �t��4̮n���� �b"M\F1J�	I(��Nhe�I��b*;�3)"L0#�Фt�e[S;��N���3�NB���*/�_V��ԈYw���[6�[�J}5�+D?�L�ٝB��O�'�Ki3��R��fǾ��:k���K�=��sw�M��^��dE�֍�$:ֻ F"�xz�R������	="�D+C����\8����`��`�[y�8�r����i=6ٶU�R�@�O�+u��z�A�w&@�x�eSuKh�m�^~h��;�5�oOH�ۗk��Q������I�?�S�#�)�f��fq|�):�z�T2�h���O��p;�H<��Ac�ŋȍe�0<M�wYg"(�Q�<cQ���^gh�Z��1�_.!-y"yJ9�O.(���]�#gE�6����~a�og��q}M�k�-�)�m[Y�Ȓ�`N̏����B���s9�/�e��RK�_���'5~�w�4�Ư����?Op��~�=��QVf�oDs��.�I��nQ���i{�'+�Ԝ!xmŧ�<�%m/{ML�H.ʔ1g�8�Pz}�9̅\��hFw%]��k��Ӷ��ɝ�w�=�}@��m���=�.��g�����ؒ�9�nQ@�(��ݦv���ҹޘW_;��;J��F�� *�	��N����u���'yX��Y�,�G累�#��g_�
�U/�y�A&��c`A=m��v��.Ӡ9���6�E=p�v�zyz�����Ք$�94�=^^�y��BۯJHiU�9����q�0�Ϝ&6���oaύr������H��bim��6�ljs��À%X�l?�,G�{䍒�Sd�ܼ��V����I�']OQ�Z8)��09��<&�3i�߯'^���������nf�R.Ў�K��k}����Q�2��RnWEl*��eN�D��!o���CQPlp���%^ؿ��p�S���ϋ�N"�0X�:�� }p�yN���aړ't�4B͑8��-����X?e2���i�G�F�I\XƯ�����\��|����Z�ٞ?�O����:H��Y/�j �{���j�n��~FE]v����^v������~���!�p�NhӄwZZ��v(!*��,��c{���1<�c�	�>J-���k�յ,��$4Oj�ǅ7��)�c[3�B��G����!������KIj�ƍ8�����G�^Ί�ߊ�M^�oq�
?L��ߧ�p:G�xΣ�we�^���΀��%����FQ,�P
����EC R�&.ܷ��LH[w!�&W���(;ԗo����f�ZK�8��O�C���&�k����yP*_f4�Z?�KO�--n<X��m&k!�EƮFㄫ��1�F�oP���ib���@��-;�x>cy3�\I��e12�`�Fn5>�8hg�by]�34e����ӿ ���ee��dR�y@��Dx�A1�eƎq��ن��'��2i^N̠��kt�g?�A}aܙ>t{Ou}��撉�C��&������@�� �h2� ^�Y�8܌���3��Hr��>:�,����K�ඖ9�������n��0�ᰐ���z�w*�G����zk��|����D
h�l��3N����m��K���f0��S�����k�3Xƴ^{�9'�<��}��Q�mP�;��Bc���;���_	#-
��Pz��b!4ϮI?����R2�M��*b�s���Xo�JŒ����w��O7��m*��9ߓphY��s��eA�WhFl�m�sd�A��a��d6�9�-�r���YEA�������,��"k�e`�7�S�Ro�<,(���	�r��C ���j�v���1\�,�����FC��!���lD������9��Ŏ Y����o�̕�m�����"yΦ�bn@Af�fj0�t����f���`���Ϸ���C�S���@��A�h��SH՝���jԱjl�2(������������臛�����_�4�1C�Y��Л�S.`(2�am׌,��.��Y�]vhQսޖ*�}g�}�0�F��ܽ�(��+t