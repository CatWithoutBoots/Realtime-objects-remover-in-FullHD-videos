��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�P�:Y��g����N^n�O�}G�4�0tG�"p��[.n;a^���H�jٖ��B&���$RI��d[�iX�շn5�6L�Ŋ�Tk ��ezJU��A;��2� �fg���ȹ����NK�"�&�0q�:sx�{��u��\���8|��J۫P݃x���0�F��jj�ڕw��M�|%�tn���B��N�T��<8	�Uz���j|��;�I)U��'>�@��|Ȳ�������B�c���5<�^�%I�4��5W�L�{��ʛ�;[���p��j���$���7H�PU[W��l:�ƍb�n??���'�v�oܑ���2����� �Mj��C4�,���o�2�Nfi�-���'�"��D��57~PO��/��ݐ�6l
^8w4 �/��7�0�4z�\`ƔB��=�1ԗt}"=���^ ��b״
*F�z�퀆�L	��al��t,v
��B�3m�|<툿�^y8�}%_�[?�04e�+ْ�(J��xE,a%9[%��;��5ܙ�V_,gǑҖ�"�3b���>�L:q����q A�-o=b�* �;��T���=s*�"���w�!���c-˾]�c'��o5Q�wI�^_�͔|l8w��5v�DE?ΐ�P�
���
��7��0!O70���$�J�'��ԝ;�������`LY���U8O���stK�8��F�y��
T��g_!���cl/|)�֗o�$	f��r?�G�lDw����?�q�5K<�G�;t��r�鏩Mw�t�\?�_쏗�`�J�Ddf]y�{��|�'w�ؤ �V#!͹�A�;���r��Kl�H��LU=#.�=�G�5_��hX�Ⱦ��<�?;1�F�C��+)�>��'[֋�]�qk����w�Ɏu�y��pX{��J/s>��|yj8�hICW���r@3;_9�/�ȦC��1�ZP��@'�#����N D!�J�,��O��5����!l\m� Wt2���I�B�w�?~7�=��@�GFO�9�b
�	�m��<��>V9�L�1Z�#L/i�͡H��PN �p���5
�i��3�Q�p����]"SR/b�́�Ղ]/���c����n��D���Wo�j��g�D����-�c��Թaꭄ�P��]o�1�#rRrD������Z�#g},��f��Iqyp��{ɏc����/6�ɣ��(�ih
�>����J�b!�BC�;/画�Z��m�ݖ�����7XF��+̲fG��:TgB��AQÔ��ᔤ�9+�nb�;&w
�c��8���]k��+�Ԃ����3Ԝ�P�"#�:`rx��|�I��a�)t`�$[����Ay��3�N����_T/�"�i��m$�J�qC�y@�?<���1�X���8�����lQ���`���t�Z  jEo��M��\̬�z�ٖ^:	��E:���/7j�x��\�,ɘ�c����lD�R1��`�w��ê�6�g�̚2lk����+�u<[�Q+4 X㨚�˅al���L�{J18J�n�6ּ������=K!1�n����s��1�Jl>��uFjt���K�d�\�Y{�sʴr5[5�{l3��pذ��vgS��݌��B�8�B�u�C_�ś�	PNRM �U~�̟�"�W/��6��W�fՋ��{b��%�j������&���̎9R��A�:P���l.X� �~:{�Ôx�򴵥1�t����,QŋS� O��;����ѹl3��a�_�P4d����p{�����Hao��wQ2V
�8�z�2�E���=���D��k�35�'G6��y
��9$�e�?���P�B�?9�7Cfл-�Q���y<��Ug7~'u�R�-WY��~X� �\�ɢKo�����!�:i'v{݇�N��c��"�Y� ���!��b���Å�R�Y���4��0��ÛU���鶂�t6&y4-Q7F�f�ۜc�py��oԦ� q?����e
~+�f@�����T-���p���5�\�\^p���'X� �>��v��٪�R��������c��+\����{"���6���dH�����r�fCȔ�����2"���;^�f��x��	RK�_��Z��[�p�ρ�n��0�{��G�*�����
O�y�"b-~�'�/�
I�K|R�W��T&M��^F�}�vk�\u����@)nK�zF�T0�ue��X��V��i+��HT�c������|F�߼��iȴ�K���ߡ�s��>�ܞ���C��x�׮�+鼖���=�m�����_n��c��w�H��<�RK+ce���z��'%�w���0O�d-*�a т�4\�<f���L��T~�?
U��*�xuF��a����HV��{`m��}���'�L4��i��S6r~��3"����4پ\t ��g���&L���;�~�������������8�!c�ǩL����̖ؔ���>K�uz�7M���SF��q�ϣJ&'r&�7PR��p�\�m��i�a�,�7�ľl�dq~Wؚk����&��"��� ڊ+��y>C������&���یa��[�a*k@�@���6ζke��=��۰��Yi�����V�e��`�[�H���RV7�z�=8��3�z�{�2B��p:��ive%D,&���������&�FڥB��� >�gE+��B]�.?�	�in��#���'�"Ԣj�@e>�#��t�>�?�h��R��ƻzI��DR�5��� ��1�)�-�5�,��K:ET���0�ݠ��Ǜh��&�ÄA]����i}8)bo������"�ot-zb
N��({5���dL=�Qc��~yC'�:�tGؽ5y����f�j�G��F��$�đF)��{�Z�ުƳ��&���9��'�"��H�X�H5bI´�h��?�^t�#q��gC���k�#�3#���E��s�w�]���bJ��}�': t�� '��,�/M1�G�ͺY���hFS�?�nÃmV�$7.{3m�#��b��ۏ�!�1�%�� Ø�3�.��$@J%#�5P_s�y��HC�m<�()���74���<�"O�-�2S�F5��q�x�q�Fl�%ԡA�6>���+�JBXD:ac���,��d3�]na���BA�E�(B�C����1-z�`��ָ_��%*_?n4��Ƚ\��7t��#j��]Ø�#I� 8 ?^f]�I�|�E��H�-Vq��<]
��0���գM|��T"��#r!���bP����0�Nr��P�a����H��A��ͼ�g�"5�#�4A�H�@��Cl�/D	~A���Vێ!;�{��=�Zˉ?��b�:��
'sy�P)�ħ�͒N5�m�:u	���ː�[��,"W)�"HXҳ)�#ԩic �+,\�{�V��sS�W>����f�X?B��p��19�=)�1�,).��a���G5.������H<*ɋ��L���/�,��0v�M\jM�2�5�����_�ςe�J�TNZmJi�� �JC�'RO|��Ki�B�F�� ���u/.9
	��d�#V <o!��-��
G<Đ8o����p������3�g����K��]u�|Q�� v��lΰ���L��Q��|T�3��(��Aܧ��;�Kva(Y>����b�v")�C�A��v��a���Y��f��)j!�E��_���8�����H�`!��d�f��@��7y4�w3��2<ė��e�Xx�`�=Ǫ v���K�0���-��%��7Az�|���)������S����$�dw���
���<�*"k��CC�aԿ�Ɔ��31������d9�-�&�����tU��Z��H!�G\��ʯ�t�>�b��Y�
�)�����B�q��r��ôv�[:����ـ�
Mc������!�;�����`q���H�p��1�ܬ���k��,z�$j���2O�<�i�ZY-��zQ\?0�3����~V9,Rc�g��Aq�w�(7ˊQ�
��ʺ���u�J�IN�K�8:g�Kp��LZM6Z���j�$�'�8�BO|���Q�܍ws�BX�`ɏ�{�I�R1M���؋޹q��L���k�N�i�
��X{^�yy+^�	�����@_�ak ����Z�S௻��5ﾙ�X*!�.��FڭW��Z��w!���be>5x��d��1y��Q�/��@��n��"���'h�s�Ȍ�'|�!=&KR�+�C��=��
��`S��
Q>5�Ño�(�3?�4�Q�+0����8t����D�!�~�6��?�>�|1��c����{���B�#RC�J�T~[�m�^ۉS�L�v��ٮ#��0_g�m�#8�T=F������<P��V����q��L��c1hj��ŗ�.�����z5(ү�J��f�j3R/Ҹ��O�׫E�"�̳�	�ɲ`W�m@d���A%�
>��X��1�S]F-�2��e{rŝ�t�_���%yS�B���~
PG��/��lfR��6��]�f�`J�Z�����X����"�ԒQBzmc|���f���.���<�)�#���zDP�˪z@���bR5�$4C��Jlrb�6VTI����+!9GƱt��Ϩx0}���j���l\�����u圙�& �6����1u ����A���^����ya�V��X|���K/��@鬟�< �v�`W���,PL��0���IPj�W��0��+�ئ�K0�C��CW��}���il���<�ѷ�㤐�H�aX���>� ��$��v��ԋ'�*��-	r���^��F3�W	
�>φ^^z�	�4]���9�R��&\�94ǿ��R��8tU&n��ʩ�>m]l��{��;���B��j�'�v��~����j�.b�%��y?}.��ỻqP�q��XT΋��]2�G�/�G.B��>P�X��W���5?G���27� �h���0:�D���6�2GvM�=z� a(Ēy��ǋ؄��Z��,�#���и�����V
�_W�AK�Z�3��n﵉\���sNE����^ל����� J��!@�	c��Z8Bf���&<��i�A�
<��q�����&ǃ �T�G`�yd����P���ĸ�-i �+�t����Kt�l�p'P��CiL.���V����&N�����b;���w&���a�9���"�J�1��v��b7pG3f���	�M2ò��5�ؼa�?���Ȉp�,r ~��:����7�y����f"R�E���'��S%]�mA��da�
������8�%�?��1���,��C����r}ㄽJ���"��
�Dǿ(���BAkɝJޢӟ��$���6����k9����il���V�6�s*;��/���G��$p0Rn��]��*�/Ɵ��\8H=/��49��"v$Jד搦�C; �J�a��!H�c�g�ԈJ��O��3?���R�W�R^G�s�J���cPG����.����khvi=ӾT�ě�;^[d2��+��ž���?M��~1��ӌ���'��U�iՂ��Au}f��%.\�����C��h��T� ?�ze�=���g�K�n�,i�j�����m�Gc���$�[��V����UK�B<�('tu�4O-�w"Ѷ�.'5����v�Uk��~�����	@���hr'������t��[}LU&X��*��b
d"�6ĝ�Nُߏ���b
cf2��ģf�h�"d�������yIƉ�xNi" {�d��RZ5x�3�us����(����>a�׵���3��B�o���\�k�9�$���߬�=։���P3C,C�02M�{��Y)�!7!���3���g#w #B���$[Ѷ��c��-�zl:.�Z#J�E &�.�u�I�yX��B�Y���jI] 9�T�)�յ5�Y�)g{�ugj��q.���^L��k#�'W�p�<J>�T�7��h��լ�r.T��u�����}��,/��".��N)5�Ni��΍_�?��\T2�wetH���o}h1��r���r)N&�xy�d�D��%��g�����NY�Q7�S�f~�h˨��X�;hOy����'q�<<o<>�Ss��}�	��x0�/���^��:;�|-&z�U�MM,���d'%
rH�ъ̈́ 6�]�l���|Si������J�E���O�肆�P���L�h��c�#�������I��QJp=E><#'�)1$��[���~|�S�������BƟ�H�Lj������z�ߚQ@I�+����+��e��a.4z�!Xa�y������9�h:�{c0S���mZ+�9,����'������l�?��$��c�n����C%#/��LJʯ~��=��׹����Oi��[��7�;6~���Ҍ�]�U�#D��$�(EK�wB��%u���W��b���^V5a�|�B�*��u='$��s���Z�i����mq��7�͕0���&e�O���w�Ws��,=&>mh�+tWrL���\r@����W��A��7��?q�j-m�
}r�:6ޛ�i��C���Y�S��*'���2	y��-]+�mm������FB��$���."&����'(6�j�\��!�QJf�S����>��aS�ϲ��E�>*V�.��������mh�ȵD�Y�n{0�u*0�}4���F;�V�Iد}C�q�5j ���{��K���3���׶ߥ�B��\<�KL�rڌq�>a��`��,Z�����i�7d�o�Ⱦ�-����]ZJ����=�RJ����/"�ob�о��J\sR#8�.<�� �%9I��O����|X�Q�D��Y���y~ ���:Cp ���f�Ζ��m+�X�#����� q ���Xko��{��n�)�c6���LU�/�{2M^l�p��`'�:���x�����F�}��V��V���b�p�b/H=B�� �/C����ף�]�f����E� J;�I�o���Pt�lbb�
<���y^!��У�p�-��QjJ����l�Q�(�z��>o�&h�]y;�������Nh�$�	!o�%%�_$�F�z����������C�O���֯�A]��v�( �݌��[��h�ɏ���0K�fV����<��BİZ��3	�\2d�kkBcCc�ܖ,)7JWw��i���|��� ��0=�	��yn:\�7-V_����.�پ��^1L�����b@�T u����	�*b��+�m0Ym��#Pp��df���lS�ļ��'���J�����lzsW��xyƈb������k1Q� �N󫆋�i�L*g�/9�?Z�/S1��+�)��&�0�F��v�<�>)�~�G@6R�|�]�*1C;�+^'�Z��h��e�|#4~��y�l@1"���>76<?�e���̻3	�\