��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&�\a��YV4����Rj*�n��4oM��>������ɾ%�n`�*+�� ��A1�h�b�Ф����a΍���d�ԁ	#���}�K��T���aS�mux�O^@_$V��ݬI��l�&`M7qG����a��"�����:��-��WM��T������`s�C�Ҋ�,؅��n��pc��w���Kj�/��j�O)��&hPW51�[����\o��,A1*�x�pxA�.�L�	��R)il|́����=ߘ�`��{n�s;����[n��N�1�V|m���	��;O�t�l؆W_M�_�f�
qo"�e�b�PF���e�|X��-�0|��d�|�\��O	%���{���+�=%�؀�ы�Y�j�L��TA+��V���D�۞��Cm��|9�B&�g�2���F��dAo�*f$#z��yn�4���Z���%���>b�:�vo-���d��B_��т��@2S�O��&h2���S��J�3zF��7�(�R�NYN��aqM��YE�P[���_=3W"�|����ZW��/G��$>�9-iN|�j��ݓ�Y_�z��0m�ߜ���)���:�#T��g�)�@���p�}�}����F�k�$�`ug�?c��&�4�Ws
b�2o0����x�Ts�%�5��R$�&*��������@{��u�u����'�gk�VF����I�T B�4�tK�q�}�����g`�*.�[�iM=�Z<�J�C�����ƿ�յ���o�'L��F���>�`��[���UD��>M�bF���ħ�W�7�pG�O�-������$�2	\�����$ϩ����p��cק\��CD>�H�,Q���"Du��ᙅ�yG�P��%[�W���t���ӕ^N*������
A�����/<��#Ux0V���"�H��+�2l��h��v̶�4%zS0Q��kcۣ��,#T��1��8=�{�y����xq�Q}c�IƇ���tZ���� x=�A��/�f�q�CtM;i*����ߎ�{3�Ј��.��+��qf�4^�A�׸���ģRY>	���7P��}/�}�\�s�>Ը�((�x��DY+Ѵ��$@�:��u��כ�MX�OW6u)�+�1Xvf�+�n<� e�}w�:H�ԏob���CW��ؖ�{��wμ�428��
=�zh��x������������SK&5W�+&r|�i��xć�
zC\&L��~���%���K2 p0C%>���P�"6빠~e�ed��J�4�1��\��l�B�#��a�)A%~�&8?�e��N�h��\ߐۛ�������1�h����/�J��*�5�B��T
���|�&�rGK!g��ݝK8�Q����_��H��S����F���v�g���@	��wwJQ�3�KK���C���Y�s�!%���(Y	n�S�<����ą��?�E�b����F�����Á�K��4����<k����㹂z���-�zP� ����]?�'�x%mpv�`c6�8��3>�W�;��k��y���A6��j�Y���@�[�[/���⾅y��
� %����ӞP%�LN�oy(�a+6b(3Ϥ�m,���<`�*�q��[:�]ruaϯW���]_���	���L	R-�@s3��ZU��K�1y�[�&�0��$���y��:�:D��fO�`���r�E�����L��WQ[�V�FI�������P�U���AN$�/�b^���X���=��m���ſХ;!LG�=���S|W�+1��A�X��2,� ��2G���[�c��~�l HV����}����$�t����uJG�s�9���0/^�yQ�QtO.M]^�sH����t7� ��/#_��)VV3�_
�ئv�Zg1p0ɹ�Y�L�F�s���ϲ�:��#�j$^}ڳ��^��̃\��wg.�A�-��#�>�'(�g�Ӟ�M��І�(�5�S���9U��W�rϥKx���x��A�Q�!u*���� �3Y�zl�KR�\�
�^,�Ȇ?�`P���(�rؙZ�@�C���Ds�/�Aa�*�](�p�Ѽ�b`Н��x-����e?PY�F�ХI`��b2��{w?��Ҿg-��[���R����|O0_��8���.D�+t�N�o�Q���������B[���*�o���%��n��%�_�Ȝ}3�����sn��F�|�M�O\����Zhn��dj2�|g��X�D;j�<&;�:shl3/�,Z��y��M>y��<�i�2]��@_
�����07�I�l��`���h�DCc>�[����6tC;Lg�>�l��Z���h8t������h��+��[�[L.~���0n��}`��K�*������i��bbIB�������l=�o���ʘ{�E�N�y%��b�-�n':��~�����Ur���E)ݦ��<UgpheX�-��ɪ�B'������=�T�M[�wuL��Q�H��@��/�BO�)C�:C�
g�:�"�׫k�.A���ac���)Ŷ�
�$!�n�4��>L�ki�b-���S+��-;	fi?�lQ)"�����՗�P���m{u|p�Ԗ��p�ĸ|�Jy�K��m�?ob H)���O;�5�\��D���@��{E����g���L�z;5:O�.�^��Y��8�!RqJ.��W 6��
j4W��!V�JEɽr����.'�cY�}r�I��<��r)����r]������$X�|��.���I�Y ��|#����l��i��s��h�!�v��d<."��L��}��LTrZjf�.����⍠��aF	d�q���7��������cwf=�J�3<���':�Q�뜟�scc���*�(�A����4cj��~�&T�?q�d`��̺��ҟv�Q���2�y�E���U�+Ă�l͞-wK%��¡%~=K6��w\?���$_��j��EDUӦ:������S��Dx���h��P��fwP2���]s����X#tV�ي��s�y�ג�};G�v+�#+���U9��~����(G�V��jݦ�O�S"PA� � `7��X.5����| �d��O{�&[��,h>_4�k�=k����X��/��+��J7��<'��t�����C#ETKs�ԙ�w��o��"6�kje�f{𐋺�ɒ��n׼�W�H����+���!̳9�?��-����#�to2Jz��ϛ�]7�΁
��.�������Q�~[�0�3}Fe�0�vX`~�3�aF&����)sW�J�*�jP� h�d�O�l�]�`�w᫇ZE�&:F�ln}�!h��!�80q�kb%�d߫|�)�9�8���.��>�]�9,��Y@�6x��5Vor�C�mBF&	�r�Jv�۰'�H�t�9Z�������Z��!э�`�a*\���(����Ƣ�w��j����tp��%|/�k���cg����C���5�oʕ5f�I���!=���E�����P�J	�;��H9$��)�K�3�&���C�C��"]ʸ�N�F�z
�.����cc�4�	�a��*��ks涛3k���'!�:KGՁs�P�v��g��M�~v�a5���(�/r�Bc�(+Z�)W������ꉲ��⿝�3"������m�%^F$����~��e��pS0�Qm�O�a�sq������'�Ճ�2�,}�Cvs(͑�aV������5���{�j��3�#�7
6�MM���π��[�㛼/>�E?:�o������ �vɘ8ܳs���ȴ�K��)Tz��1yy������pQ����@l��(d�`�w��ɹ7� p@^0-�k�J��wy�D=� `E	��c`�­�.A1��#T���5EH�1$�`Pw����e����t\�4��:e$`W��s%��?5	T��'0�k.9�s�5�r^��/b�\���?��M�K�����+�P�;f	ɼ�٦�B��Қ0��,�����;f5Xw�ln� �v.] I�k��Fi��D���<]���O��"ʰKqޟe�"n&�;�+RI����x��;~%�A疬�ьrth���N�Jʨ�t~��T��v�θ6�����#���:��L��u�5m��2=}?��ٓ
G�$Z�)#KVH捬B�}3�jp��s�B_����q��b��#K*�|�6��x<_��]Rn�a�xBھ�5p�|�����ڃ�g�d<h�R���236�?^�4Q�i��by)�u-F�P����d�`���bǃ.6�����-�,Ў����l��:~���Z.�9L�ڵ��:һ/�9��y�s����f�1x�07<sql���0��%�7�t}��Th&��#��Z�⌾y��E��
��g�'��ܲW��ם�镗�ۀ2�����~�n�Hr�t���rdH�J�$ ��^�Zz0C૫;�d� I�,�Ϧ�ça���n3�| $l:1|o�����	���+��5���HLOQ�7�h�K˳-M?0cR�%v �K�Rw�����]�J�Nb���lG����\�5�[�t=םd��_�������b����	�ό��ڇ=7^��a�����/u�`�w/j.f�7c)p��~wb��������A��I���a��w��f�*��6��C4��߿���Y��_�ϻR�ٰ �RZ4�P�46v��-�4N�{��C��Bu�1��w;��d�@������D�V�]jf��tU��k�4vx��w�X���.� g��	qΙH�+'��H�l����B[m�j��\�D�����K�b��6p�uh}�R�(-�wa}h��m���9���*�ȡ�bj�׳<��~����ct(��J,�L�<���>�r<�`��H��� ��u�?����,}���F�0l��߁D�ED��e+�ȷ�&�Cs*��:�P�խ���BD�˓�𿠢a+���%�0/v�:PѴ�P&1};v����>{ơ����|Qs$���`Q���Ơp��t���y �H��UXj�ʥ�DӺWeS��6�SX�$��u��Ye�������.9尙�b�)��: ���V"V���B��gĂiy`d`' ,�(?�����R`��X�~l�P�O��Y�&SG��ٗP׏�-W�,��)�8
�b�3� qa�Z��[�~Ԭ��cu��j������Y��i�e�D�f���5��1�q�3��7�)q�H�#�FNMj����F���x�
?�����a�Q���GD8���dc�z��ow�O�V�^JZ�59��ZG���y(����\�+��n��晑]��W ��8'QD��C[*�����o��&�y�O���G�za='J���ɴw�f�uo�s!B��Z)��8���(�7Q�KG7jSN�˶roT�V��LA2�3��+w��d�9b��-q�Yi���a��o�9/�3U5�w1A��bTצ��3>�.�����Ֆ@��.Մ����5{���E=�a,k �`0;�#ų�3�a͠�����8���eR�
O1�ݰ��'ی˫nC�l�(���Σ�h��)��Ж%k��$��đ��"N�(5c���T �B���$Q��bN��sH�a�{��x�R爜�SxD\�N��ԟB��|
�+i`���c�F*;K�E�<��-���]�w�����8�^���ype���A@�"%5�M����L,�H���i��(�giج/|X�-8��O��#��C���S�:N��y��nC��	g3��e��D�;=�7����&�ܢTkH�֔jR�	]��q�}�bq��
@�	��xZ����Ak���:.�#���	�ꏩ.�Њ�d�}�Ͻ�Ŏ�ˢ�,������=�T��.��s�!zL��Z�8A�H�!�h(38{�1g져L�ɟU6��������&v�_�����-%��e/�O�����bj���+��|�|V�Zᑁ������_�@Ai=D�M[�����p��S<�����L��JW�T�B�)H+�ʦ\"���Q7B7X�J���.i��)FF]Vf����>��+���� �&���Oc��609o�V�Q?0�پ��U���k������v?�K(*4�� ������H�9x�A�R˃���UÙAݩG���$^��4�ɸ�A̙W���t�˷6LfO���;��̓��杍n�1��6��U1\�~��*t��}�]�
gK�
�����c҃q�&��ѐ�mq�Bx&#�dҦ�!�I�?����(�!7�ӛ#U�H���� ̌��$0�V9��P����A������;��JaM�7ﭞ5JL�����\2.p�	餯���>�����q�k���_��o ����'��(�=�ѭu6�$Qd��� ��Y�����z<o1}��h�z`Vc�ŌɈ�.7L�r6I��RJh=��e�qDL�%7z{��*��b�\�.,���#/d�5B*��_�����(�D3���2�D��V,�yXN�:vu����sh��y-�|nt�r)!��K�p+p�v*��Ĩ&�՘��#D��?/�	���nl��7�\�V�<�-�)9��'���b �z|600����\�}�"p' �.����4��Tˁ;_i�*��=�?�����b~`�&�tj
�,h�G|�D	��_K�l��Cf�>���h��O�����	�'��;��o��Z���)�V9�R��w�12�G�#����fɱik"���g����/� iF�6�`$n�5"q����$��]#��\ �Z������ɩ��~}Ȍ�6���I
:��ݟ�&	��Cp�{��$������-�/0Y[��gcbܱ���L	��yܻ�����8B�b&�T+U��Dp�>���R�*V+ޜ�A��V��-#��"ku��.<��pB������/k��'��'-� ʎ�T'Q�.��e�����J��H-����%���]D��:��� 	�Z�ƙ��F&��Ќ�Mcb��O�䄕%=����	����z:�X-����J�>Qb�;��M��7�8"�R�G������4�?]����	������'���,�z��o�B��j��۸����D9֢�O�7F/`J����2�K��]:V;�����.���s�S�m��硎UP�����v�WT&f�o��bh��o^�Kv��ZE�~�u�w1� �:u���d(G�kU�K�Mˡ��!�v����n��*Z�q�m��ލ�[ܯ�g8���h�+�
1g�5����cڈ�܍7�fgN��ϱ�$@�w�fZNߴ�`�����{��b�@�S%A�f�sv���g��:��0j�����(��)X���h�e.�@Bs�<P�(�T����E�b�a�	����7j����ZO�]�^
��5eFv@��D樹��d�%���'sը��
H�kM�ȑ�]ŉ�<X�n�8��&&UA9|�Ə�����O�F���ҙ��%6�Ȁ���|���v}L7����9�u�S4��_Y@vFUe�����8M��ˢ��9zS�Cn;9>~w�J���X�?�¨��C�������x?V\���G��W�ƱT2X���ۙY_۾z�h&��w�g/Ռ0MT&�������l��W�eJ��H�d����rv���^R��bE��7] �$܅g���wY-���܍^�� ��\ȵoщ�,!':�����j�G� Z��C�-��|_���JG&�xҩSZıtN�����%���h����]�X�؈���^�"�.�`���2�=��Z`�ea,3ZAX���xG�F�a�|/H�A=7Y��X���#��:��A8b�&���w��R�C��y�;�m�mJp���7Tz9*�r��P�%�A��;{��%�@/Fy��{k�ĐcZf�ͭ�2����Y���	��>�X��Sdgօ������y�����=<W�w�������|q}հȶ��Kҗ��5���%�Z�1�e��	������k��Qء.�6~��ƅ`h��8,��@��l-���Y�b�E���x�2I.�x���3�!�'�!.i�ld��?x�(]
f����J.�ⅺ��� yM�y8!��:&�m9\�Dmh�ЅN�W)��Z�?��P�{��D(!�_<�c.����^�"�Dz!�>��).�-�t�x�F >uZ�	;�hF>ȖѴ�!���҇˲�Fеp�-�O'\�	��_�j�Q�FD/��M���F���1C�䇯O�����_7�zo�������-d�-�K�/�hf#4�+l<�����Y�y�?+i�[�q����F3߸V�P[���& W���+(G�v�o��
]�^d̠҇�a��/_�c�c����F�]�d�wI)�����6/�����M�&�/a�[������v]Wu��X���P��+ߗ�M�D��ܩ���ڄs�9@��N�&�FT� 3�}G3��8zQ����9�|Yr�ա�pW]n	g��=mri��Y1�< ��_J�v��!���G:��*1rtYI��3���V=��M^�,$��)��a]�w)q쮺E�Wtm�M>���J�{�E�����qSF�|�N�nΦK7PD���n��z�p���m�&�UlG^ �P丞�u�q�^'�^mCUp��J(�(k���XΠo��̐+Ā���K�,Y9V﫸��59�}��f�f]���V�gA�)���)�Ta��Ø����w��,��ܴ�o�m����Vв��B9��~Z�LLb��� $�G��;G����a���g�y��#�ت�z��oCp��=gF%sR���M=��=��Ir� 4!x�
��X�=�~�E�����|�V����ODH,2�
���e��F\���jK�;�=�[��
p7�\����9�G霿ވ��ʦ("� '�:�1ɿx���j��pa)-x!�Z%��Mm'����&�je]�����f|J'(W�d�a9��^$O�l޿�ٵҽ��>�do��� ��o}ξ���0�f��Z���x��c�Ne�'E�?�b ����/�Qoزv����[�!,<O�\7�<�S?y5.���8��`*�8&�S�@].V�B�"T��8?>��}*�G�b�L�Q��֨1+���Ҭ=��o�	ţ�����~TYz>��M�n:v����`�����y����gYR�u��H[�|TEM���e/+[Q�(�e�_�nu��T�:��[T���|E�� E阛����+�n�2K�T�"Xե��R�1���s��,�m�F;��Z�PH�2'�O��*� L��S%z�,u|;2r��Sȇ��*;{`!7^��,�1��L�ܽ�6�M#@��o�J s��$��A:n��o.۽��˻�5;�G2�J$V]Y�Ɯ����_�pd�0��	*�wmU�ga�,��(��u}���z�{��!ٷ�&���{x+���]d��H94����\���زS~�bvc��?��K�ÚX� �����Xm1U.��%�\��T	=������k6�z�qĽ��S�������W��n�9S���(�[ɟ�cp7=3_�҈���V_�Љ2�٣�n�
x��/J��8�1BȘ,�2`(��#Ne#��g p���Y�g���#��<KUT���\-�!w3�~v\߹b�,�~"ӕ ���E��(w̪�Ng^C�LS�#e�;퍬�ۦq�*�3��GA���s�[��ؠ����Lv
KM)�:����e�"ÚP��`O�F��T�()�j�(��j��ܴ������<�ԵJ��̻�R��L�)�z���c�u�8��ے6�ڇ���1QG�X'����UΣ	[�5�`KW��Ra<b36�4E۰��͐_}��{C�|M|H5�Qԉ̱*�ɐ�(�r��{��?W}����G��:��csf%���Yt�4�&�+)G=)��_86"�������L�w��%v��`M	�������u�S�~*�˄*B�[-,}�^U���ws,76 J~���++=��!�ԫ	N�w4����g<��7*��z���&�B��.���n,��0���ߏ����!�\��ox+4v���1_�X�?Mz:� "����Q\� n�|��/S�a9�#EҠ4���aMT"�coB!qB2j������k�#�4�S�WpyE��A����~AK��UЅ�o���[&�e���S�H�	��|ta�����<�b]�	��:�����1^O��L5���ꏼ��?ؿ7���(��TSR��|�A�Z�}?ɰ<{á��R�Q�]�4ڟ���UL����Y�u̑TW�i��jf��to���ԝ�q9nΗi;!�d�}c�q<l�cߠWb�I��{{4K�mm���<yR��Vo�>�Yn�W��$Oa�+�%5 �Vr�e�Ud\��R���#sw�b�ȷ0��$�W<@f��v��0����C'֌�A#M���ܘZ�g(n�o���"��K���A��n�$������dX��aĴ�� �7?�6�&���k��
��o���*���F�D��׆��)/��Q׵JDDj�]��{e�s���I&���aJ�gw�}���F�lrC�����
 ��������|��2q��z31�����Ra�y�_�U�.^SJ���Gg����` ��X3� �e��Ol����&�(2#�Y�0r��Xm �P�W�e��-����6��េ�����|r�.9��r#RD��hz�`O����ܞl�므v9|u�IH��8uZ��	%���R�Y�$��j6��:��jJ���j7�}��J�����ǿFÐ)��Z�AV���=�>:"������(�� GH�p�4�L�N��"jn��c��E����K����4u�w��9Ȋ�0B-;o�D1y}���>/�����Ŗ�X	�[� ��*����
Q����ɘ3�Ɍ���x���2e薡w�K�H>o����+j!�P�t�k���݉���f˜��X���-�y���в��4��I�X� t�0Q��;J�.XJ�R��:_��	I�=Ы>'���	���+��2H��DM�Ԯ�@Tj��.5�����{�����]���?p_xy�?ʊ��߅�oN�"��6n�D�4����^��
��J.Ѐu�ǖ�+��O����f��Y,�E��㱀��Z*�VP,�}�K(���|��D�
?�p<;������^�[%�4�J�vwKRx��!�&��ߺ�H,�s�ٔ�'��b��w,X��IX<�}�-��ە�Tڮ�6j�k��A�� ��n>����$�|��-u�|R�	����`��Z��	i�H�n�ԯ)57Y��&6x�b[m�����X��g��鹚��S�:��d^��g��6�l���k��=���=��vr���uR��&�$9j�[�K��8.�i��\��Ț)![���Fk�]x����2�ݿcPo�F���*�&�J�Mt��A�K5=�yR�8qd�S���j;F#6>�?9W���6>��7)�.�����F8��ˢ��J6��|Z�M����VE��>e�x�Q�����D�UT�aW}���Ù�v{�a�n�||mv:�E"�ri[c@ ~N����O*�t���� �[ʽ�dZ�U�08����r&���YE���.9Ԃ������ �N�:#��Lpd� �\����P\�n��HO�u�v�ktFNJO.h�����X&��'�M^C��ۊ�%��\�r�.��*��:���!�9a)]%LF��>W�	[d�~d!Z�/����X]�8�ȯ-���r�Ƣ5�����)^����u�u\��ľ�pcS�Qj%���4N��T��v�
N"O����?B��a{}�1ńsB��hY;�&[z��k�(%mPon�_߳�x��,�.{�ly��s�a�[=l�+�
M�>򣤪԰]�ĽH�xV�ÏU6kς���4�`(��q��j���t]0Ew!ޡ��8����Y��[	!X�-��s��&��,߭�˔�&�ֽ��ŀB�|��F
��PITp��C:m�#wYʑ��
���r]ck�=3hc��Kd���Z�&;�e��	�pe���6�����ۮ��z5����i!��	W��=WB cE�O��=�→����Ɏ�T�w}��W�S؉D��S�r0H�C]˲;�J�!�AIHg�w�r�ze���bQaq�<��bnckv�xVI��K+m���.�b^��~�e2���Qk��6�i)u�c��*�Q
���C�'B�{G!V��0�S)rc�-mu��|�j�����8aU��n!j�EuXݦ�-����d��)qx�{@��i��.�.A]ȫԳ�;WTjp���W����a��ጸ���]��=�'�Jɐ��hG ��'8R�R2�%�eM���Ў�x��^�	Q���~��O�n	�.�?�Gx2ׅ���	^ѥ��~���yO�#���CfkR��ȇ0HgS��\����������k囩3��_H {����&�L`F�8�/ei�w�#�⅕�ۢ�I� s�ؘ�m��T)��@I?2\-���B�#UfƄh���v.bh0�4Ϋ3��V����T~�sֻ���}2�,��j`6��gC���>���bH�P���&}%B�ۻf[X��i�H@\OYڼ1��O/��&U���N[I�����٢�:3Gק��Zf�F��yK��_�9���f#,Boy���H�u���Hڊ��N2����L��)h���KvfC3��O7�c�rq�/ө��{BlU�k�����L5�-��Hl�q���ĘP � N!�&����;�z��ĥ^�b[��>po��%����lD���:��>F�A@��̴8.��w��V�c��A)6����	[V�x2i�:��ǂ���h������!6�+~#YQ�|[R�`,Q���we�\�Ky��{�
Xg�Aw�gk�8��X�LҨQ�Q5Q`<r^�+!�%�-݃�ne��_�+D���D�߃j�@u�eN]�-�/�xz�c�}����8\��;ծ�mċ��!%fI��|+��Uc(�j�5qYh$�#���站*���(U�������BM��o�jH8�����@�}}"2��R	�n�N���,���c`@�'��ڍ��z0�<@�\w2h6�=� UQ��}�8WvB�H}���0�\6u�X\9�X�W'�iÌ�I�%�t���ѬZs�"b7��U����#�-md�+���DE�@����N�@+�$4�������!��y�¼k��I\SF��S�}�@Hi���3l_D�C��%
�p�n����o�OT����i3��&�LA��Xڭ�֤�"�^2�>�s]�/=��L#b葦��RG	��H�^��ʰL�:��|	��$�A�5������v��0D����}@3�l���ڦB��������Ą��u��։�@�0��)��MB3䗐�+��*��Y��4�*���2i�ұq��T>��yxE�^�N� ࢣS��Χ���d�'$��;�s�6̈C�t#�A�/p�����R/~����$����g�6*ޛ�C��n;gK-��>c�'�sY[�h�M#�D�n����K,���H�Ҳ4�J2�p�j���s�����>�^)�N�ݣ� ��y8�h.��ȅ��;�#�hxx���/����r�ʶ5��O�T� (��-���t��LZ�AإLnHw���A�UPԅ�W͍¢d�������ow$��w�օU�S��q�s@�wZC��V'���K�19����?�ٺFB�O�Ca�]��A$:����,2�
&7�;D\�����/�4�4]t������W����I���ЈنVnR�N�<'N���>>x\���p�1Z���M�>H97�S$�˟|�4'G��i!�4�4���rW�����2;��/}?S�/�W&��;/�&}���*��Vf�%�����'��'��e�.�5z��̘h��uq@��p�j�1�KeY�]��@�g�ȍ��B����T1��)[`<R�����KN�I�[���l 4���
���ZV��>��A�g�ݢ�8�?,�*��1�oٻ�zE_�<3����nJĪ��vL��Z�h-��.Z��F����FI�V���Ns4�;�K5����f�p�"ao�݅�F6�l-���o@�g���6<#�۽En�`�����^Ud"e#���4{nz��B*�����t9i'1S��@
/6pM(�JQ��j�	��B8�g.��jrk��k�`j�J^#�캀�޸��	J�mPiVp=�K�8����f�h@}m����?��o�}���D�?[���F� �j������α�gQ���:8��K1�~��Б��*C��	��_�� I,��bk����{_��Q
���Jl'#������Ɯ0��\"�5���"��h5�$�T��!�uy�[��w��w� �L�AӞt���p��}�A��Bnx5P��LJ7h�NL�r�AO�IѸ�V�y
͠��E/�~ҷq/M�UU[���y<�]�U�Z�l�-�W9G��27^��I�OhV����q��G����.es@X���`��G�0lĨ��;R����c{Vt{p
�r!Nf���C�]�̜�����L/�{x��
]a�6��#���%I_���
�J���j^��Q6��Kƻ�Gz�QP���eǅb��s
s���Px�mI�x����G��Y9�+�V=��V;�>�
��K�{��h��{�[������J�S�g��Ue���(���/�Fg���]���]0�wx�>⌾w&u��Hf����O@V��p/���D�Bx�n��a�%3`�b	<wlvfaV��aI�J�<��ht�s���1�����;'�6�X�P���w,=��F�%��/^Z��[9�駘ehnT����
d�\`Z�B�y ��Ԟ�m�A(��3�����=���'"�8Xf��������yfI}u��.֨��J
�f��%���Cճ��]!N��m��eSll�F^���DМA뫌e��-%�Bxf���J�l�:gv��;>mq��U*W���<��v��փ��t�]u�y[��_F������{��

v]O����;Ee*�Z�ng��bM`�-����Ź�
�I(��o��%��.ٞ8i+�=�$����n����÷X�f����*8I�79��Wݨ�=�$��%�`�<ѡ�������(HR�I��N��0[\EҤSf�fVUܼ�?�i�lг%��j��aN�h�C��6P�<TNƔ�����y�I9��&�§�V1���y9���kt=�|35�a�(*�9#�|p��?k��~���i}=���W����W�<�{��me �W����[΁tͪ��,�����������,{0��ʣ�+v�޾@�,��t[@D��ڀ�!j�0���v��,l�;��� Xcv�f�?~}_�G�k{�`�V�&&����9��+J�>é�(���3U�ۥ���4oIx&A�/1=����!�)�N"ur*�m��g�[%M+��"#��oD� ,0݂�%oih�$��� �����J�JxO�����Clz���,֟��{Q��E�`j�A �;���Nǃ���� .���/���S-\�,A�Wf�W[��_"]�x��{���@��� T,�M���p���q ����]� �!�אu�rbY�S Emw�I{=;"Yu�u�ͽc���/5A��|9 ���!.���䵀��uJ����9;ˑ� 9��_�t�D���E�!u���m)2��m
�)5��g�hJ�-d֌f�}D�ӧ=��]�b�P�F#�z�I��6��D��p�ȿ/��K�gI�g����{)��V�=[̈@`x��ð
7����y���3:9�\ O��q�v�W��\B&�h\�E+�h���b8gX��:�Ӛ9:A{�h��� �7���f0�4���^�tt�{zv���f��fk�<tD�-%sf^EgMeR ! K�!�I�Ga�x(IR�K���W�n�#[��	�!U�y/wm��*j���7��!�,��_5�7F��NP4���\ߵ�#�Y�NaB�جw�nwTܹ���Y���;���{�}R�H�y�� �-k=J�r��ނ�n�{��dF4�뜞����KL;Ǎ��#�F֪m2��]�-'q~s�O5�T9uMg[Ò�:�ͦWʈ9�b�ە3�T��p�d5Ҕ��~���4Rs�����,-���l���P����G�7�d��*�1&��ŅV?�{�sU����	�E�J뜄�Yj�)��l�C�K5wz�j��V4K����l��	�QB�3��j'2ԁr�������̿�ZE��l��B;@������nwA��������| ����Dٹ6�z������>���j!��r���Ĕ� ��.����<��Xc�[�g[�_���#�d;��9��@�H�����#�;
���[�^τ&G��r�? ˀ�2�~h{��oe-����f!�Z.�{��@xܶ�E��@
�8�t�u�N���-������}��s�)c�0�D�<i�P�M�{���&��D5��#�?��m�2U9��K�tm�*4�Ew� �X]�?�?�� O�ހ���l��I@\��_;��B��!��O�4~�_��b=���\ީ�LŹ$&�\+�&� �_����6 ��ż��4m�G�k&���5��t�wvZu_�AG�.3�q3�O���{�s��e��Rj��I�3� 0��֢�.��Z=ѶK���h �����?�^7�c̈́<��Pڡx��#wf�3�G�2�o��`�:pv��z�_�i����pk�4?�[e�h��D[%~Q�wzx�f��y
4%5Q*���Ҟ����d�~�p�#�_��m~�s`�����Z�3�l:�`�i�R�rz�b���i�����kh!]��z!P�Z�ͬ�f���e���s��#ѻ�n֔���6����S��7�v�q":��_�.�Ŀc�H���{G=��SM!X�;vP�q��̾��L̈�#-!���;���,{Ww������S�{�x`��T

� ��c�X����R\i'�o׶�&R/n?�䣗	Y���5o�g�z�4!޶�Vu����ݾ������g���F��1V��e� ����8�v��p?�Ge0�؂�80)�� �<�1���NO�e_+PN��n�vh�4��(`��Uq�Sk�~��/�Z�W�r�,��s%��ӌ�4@�V����MU��re���pO��y�~
-z��ݚI�Ha��EH�<�VBOt6����2A�i��1��T+�H�
��1�X$!��TWu�Χ��'48�n8������m����ȟ���ŝ�t T
;S����p�/ʞ����GD��39g��vMc=�׻Jrk�u���E�7�u؞	 Rs����m��^������J�H�o�ML�s���X=W���j+�T��N_�tb�v�!��J��m�y޽<,�W�/TJg����Fe�"<���V{]�sޮ݊���M��ݐ���BJV��*����Bl�./;�[+�_�#���a�u�q�g�-��v�{�3i/ݎ�#�m5��\(��ȣ_5r v��$Uʨ��c�a;\�5�M��3� ��|�j��(�����K�[�n�̀�zHm8`��E_2�"Rb���\.�?�B�g%�s3:�)⻲ ��t�ʛ5�#W��WFY�¸:�y������?���Q.a#7������u����Ip6K��⏇-izV�%Ux�k~sOzq��t�	iӬZ��;�5�+�b�/��~�[�,!?&��GΩX�B��]T���1n���æ���a�Urb��EM�������D�w+%�#�����C6�t]�*F�쩯CS�g���Eώrۘ�z���{kB��M|*����y|���T.� 
 H�#Y#QВ��w����V�U?G�ŉ|g��eCa��g���{�w�a�j���CB���g%�!�� ߴ��j#n Z�z��<tf&:�J����j���E������T4��� ����J�����n��X�E&�b"X������C���a����wt>�G�%ʪ�ͥ��~\�y�>uM�;���Y�3!�yɍ�@�U,��r4G񕓖�꾋�M�ϣs���I��l:Tg&��Q!r�����~Ĩx}�EY�,��V0��x&����pl��S(H�-�l"VY7b�7,�Y]�Me1څar�����vb��2��t����T�pq�Z��X��=� �f�����fy�e\<���o��J�OۊˑE�[K�|17�Z����h��[4��͘Z�v�����$�,���.�'H2��,b�=�W�l+��f�T���{BbF$xu���!�)�T�n{��7�[V����ۨ��믁d�`{3�&�7b%���7[�`8�K�T��:
�@�]:��g0�^xC���a��.ŽJ���^�Ɂ��5��Ej�) '~S���b�=r�d��T�b���,P�;9Z����ӥ<W�Ia�T��y�^j
(6cuk��C����kTnl5�PL-G�TյY����)���T����,�P� N}�WV'c�nN��	{48Q���� �'j�N! z����f�v���$ޣ��7�^�\�Q���*3�͑d3���������G(a��+Q$�Ն8�VH�"Mr�V�ỳ��:"����|��@Gn[10Q�i����Q��ڥ�+�ۮW�W�4O�MB���� ��@>c���U��(�zx�ޥP@ٶ��߄��+޽�[Z��u�Q]31Hf�Rh��N��:Y֟��\ifN�D�J��ۨ�c:3���ނ��?�]3�����	'���yB0���~G��X�o���1��E��qg�����)�R���#��k?g�\���F U|U|<�n�9!�P]y�-ϗ���W��0��Mm���;((�"^M;I�x�Wid j�z�*����W38�݈�3WM����|�m	���[՜b[5�����"N�p�m���i�Z�^Y��h��l�[�tB=u��'�X�-O�4^�Ǿc�r�Xb���"���y��a}:���Y�G_%��
X�0�W_Z�Y@et9�Gv���3.�v���b���^'B�ż$��ӄ��[�����֭;�Q�;�
�xP���I�s��� 3����Qb�ꆣ�{�v��l��4��D0M�0���T�<��N O���uT2�����?�Ou!h����U��<;�o�5��J+����]�n��z�!��m��m@%���ȫn�i����ȱ`gA�l;ڔ�9C��l��3�K(R2����X�L��ShL5�6b"�����ڇ�ӃM� �hl�I5U��I~�������\ NA7]����)�2��3�/!��ž�@2���H.EV�SsR�.>�]&�`�ۦ$�^X}�&���N}@~ M>[�Q���'p /_� ���e��.V��Ľ����*���e��I��ȍ��wF!����Wp��!��rz_�K�y7yf �?��)�Ϸ������������:mW��W%��(|�J:0�����c����í^1�y�)��Liz��b������5�t��{F�w���%��q�'�E�{���x�b�~��wW�2>O���X���# .��7��Y����I%hd+����`�)-NuG����\�_�?(��C*3y�rޞT9{�v�wݟT6���BC���$(�٢�_JN�@�T�e±�ϧF�?޹�9�Vd�=�]�����f�DM�[ � ��^�0�k��Wo^i����U`�
�`�G�mO����Pr�`�W	��i��(/��L����8�/�WG��J�|�hw�����j���d�Ψٮ���u��DQ�����~yж�
�ۖc9���)o��)/SH#�
�qr�n޴���l+�����uK*�B��U����S[�C�39;~2M"���XjUA5�q vgG�D��4W
�L��\�U=��K��WKn˹^�
v)0yiN૟R��$��P�Ap�f�(9 �3R��T��Tp��EDS�l�q��������z�nT�>W��63E�x�ǭ`����اY���:�5���sP���&3x�����=y�o0Y1��|+����<%��R	�F�}e[�Զar�ɾjP���n�"�t(�l�̸�d�i���_��L`�2�9 RY<%��e �d�Ѝ�QI���������c;���Z�JV%Kag��+����`!�:A"̼�5�Z��9
�n��3��.Z��Ǟ��ktt>u2���Tr^��32���&���w{�P.��g͜��N�~�H��N}��Px} z�qZ�)����1O_�Ji��#�W��Y.�9��ZW�ɧ`�c�������&_���w�J�d���u��/��ٝ�@���cv�!�
5�K�s}�S[��|G�Iۨt�]$�*|Ƌ_[�'"5�����yd`�0�.�n����&����)�87y��c����	V�����(�qkse[8 �毬GY3����x���'�
����n�^]�~��mM;FY@0�Qq��Y0��﷊b �kS<�G3�����uvH��c%�w�'�F�~9�"��ޮ��2�b��Ie��3�����TJs��wT���������)���LUY��0�v{=�䋱��U�~��������$�׵�S*�d����n��7#Л6����lP|�a:R��wF0��r��9v�bC,D�L?W��P��qt9�P�^f����èkz{�3�N�W�M��A�bk2����(�g;�	����3�.v����~¶���mBD\;����&8s�iQ[��U�%	��T���Ij*Gx|rpP���\�J���H����bw(Tk�����ǝ՞��Sd��ϕ'�����AJ�m�R�qrY��Q��(c3��i��������Bzk^V��r$�u�ƫ�9���,�V9�Od7��u�.ΐ%�]h͹t#�< �1��**������@��;��2,������햮?jm�^[�c�4�mK �iS�1x�Z��z{/HH(?�g2/��/���a�\�����1ק~��'`<<?���;�����xT�ڋ��z�-]�	f^[�2MO���
�FҁQj�s����6΀��w<*��"B�"�B�g|�y�����B�Q���u'�]E��h��Pw�#�;|x/�Yx+����c3�9�|�7`B��`�:�X���/(�f�*�ׁ��^�\`�e<Ϸ�$��N���$�;��<8�*�<�j:�B��
��E�?�h;�0�����ig�(|���<t�<��'1�f)G�[����T_)���=�iCЅ��.�nyz�HC/���3�{�|�c�S�ʷ t�=e�N��~�*6�mY-Z�U�!����V��)!�R,+��Ɍ)��0��LoU�+�c�Z�� yg�>&@��,��MK����I嵍�1�KN �]����ڗ�bˬS��.G֞:��� ���W�C^E���~�\!��'��< ��(�%�X���Q�=������Y�C�-b��G���L��"��F�ၻ��ӥ�o�@૟��!���2~1�XU���ߌ�I�g\��
zr���V�㱌�u�Ѝ����`f�x�6��T;l�\X}��}�ŤfG:o��G�_J�q������i4
nZ�Dd�:�?Y�Z��D<ɺ�i!:��8��x�q<�A{�kG4�:���WJ֠d�	�ݫ��2�w�Igri+I�@+��r�/Rа|�Yf�-��H�#���,J�(xrl��]�s��bk�	ΊN�n��L���ٵA�\-���6~�{�;y)y��|禿�9���ܧ@R�ދ���[>0Kl��+��-�0.c����w�U���.b��E���� g��&N���[�w
o�1Nz8I-����y�fͨ'�F�㓄^�2��I-�v]ע�_}��-P<�wϧ���<f������u��G	0�d� s���[�oף�A+R��x�T��L_%"�:N�x����6�f�����>���2�շ*�U:�ɷy�io�(��t�q;b�A�v_�OE_�����[A�ׂ|�\�<_W�	�4�Vp+�����T�.x)Q�3�O��Z�c�{��~�@c�\�Ѷp��?$ؓ5㢨��r�������f*j�C�+F��1'%%�l9�Y9~��D���h��3ux��Q����52O��\a�%¥��@����"�z��j��T�5������2�7~��zU���!����-�-��p/ag��^��6���$�nz�+�� �7��oqA�7��-�(Q0�`�[~?�#�M��j�d���;�ϸ_����b=��5���؟7	��U?^�pjn�M$-`��n���:~Mk���\~9��P��^9l:��س�'b���$>�g��]�{] �iFC 4�wq`��.�X����,�"t ��Tgs$�rT����c��Ň�B7�:����� ��8��eAf�"7rw�3ȅ������M2��lv�ND+�X(�CZ���;д�/c����[!F���k��\OҀfyY4�kj�а��w	�ҡ��Ԝ�F�״z@m��o�꽊�L��n��=i� "�l�:�����4�W_�$H��7���"�`Zv��7�+�5���p�K�P�Rx:�J��&�b�/u;㌍����֔�D�H5���I#+�����v?n��X
��1�M�Klr	�������|�����VE��t�����8�l���t>KY�5�8?p�a�T8�ڐsy�3���R�G����ä�f)��W��� �f�e���o�I�<��	�SUࡗ��O��'7����\ +\�E�wמ�0���9��� ܙ��f= �M�H����Z�ᶷ�o�\wZ�R7���{�+�CB���̀�����۞�,lk1!$	�`��|8��v�B��6��Ii=�?���F