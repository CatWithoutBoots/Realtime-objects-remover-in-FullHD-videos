��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&r�F���oh�hi'n�į.2�-`(��O��%z_+J�"JX9�O�/�7hU[��X&���{���A(yKn��E�7��rz���Fb��B�@Ԡ��g��
�}}m���@o�q h�M�9�rp���ȡ�"��s��L}�-��6��Q�V:��"��zUl��d��%ٻ��
�$����`ira��ƈ�*�d�Β���mk1���\[ S�~���R��u����������l��i�k�76�xqBwv�շJε�V����c�´�_��l���a	�� �Тy�J�I�h����:�Qi��76��b1��4���U���3҂�!|z��3+�!�-/H@�� ��c%�\#k#�Ĺ��`��}�Bzƭ�M|6*��
�m�=%��(���/�FsN�c�Y8���:îʔ����=@ΐ��x��[��gD��Ə3�>�	?�)����YC
K�p��|�LY{GM^l_��6Ƃ��ה���DЙ.c,�P����emhl~lX��/�՗=����)���|׮RR�W�SWe�����{�'���a�6������7�k:�����@>;%�QC�R�i�<t�rcp�l~�=C�hU��$����k�_���-�Of+ڪ��RvI*��A�^�W1܇�_cvMW١fA���XzΟq<g ��)䌦tz���~P͔�l��Q��Y9���ܧ���0���6D�N2f-n���/`Gf�����I���G��C{В�U�'Z>\�Gmޫ2%s�R|�;��2�3?[*Z^F
��?Ӎ����'�ҽa��s���zt�q�?|&Im��7��|oe�m�����󼹉EaE�F�Cu9���	���,{�F:����8^��G����(�(E��	�v��;N>�K�.��+G���@S��\֋G!�P�.J&����zH�czI\_d��wу�����a�۶�I��|'z𡠊Z^c:�J���VV��/���7��|�f�v�$���S�BQZ��
Kw�t��m�Ωn�5�`�S���$��N0眉��{6����2堗�
����4���y��O�¥�k�Σ����ϱ"b���� ߾���]/>?�(����̞�tbju��ȉ�'}p�}�eu�vye.�XmRz��iz�'����[�~�s�+��3�^8�elb�6�|�n�A��� �FP3�����R��q.�i�����uu�'I�L\��zMCve�O�ߐ��7lh�)}7H2�j�b���M�W<�`fO����V�*��d�N�b��&w����L���4���l�K�/w�w��\#j�-^�Gݼwp��bI����f�����)�U�*����n����"lW����N��j
ֶq$�օݣ�xZ�m�O��5�Q�3��s��l�bai�~��S�����qKM�M0�,k�~���x)�ixJX�.�1XU�ck����+�B|�rC���R_n�6�c�K��*�"��r �;��j��X?�8cF�ުn+��l�t�`�Q?f}�������ոC0�x0�0�(WV�.`��/��_[2��Uf���߫9mq�$�iBg�������/�-^)�[h�!H�ԫ�n�bfX��D;��`��&n}��0��y�)�_]�@���M�¾zH�[N=(x9�Z_Fu˶p�m�����s���'�9���Hp�/=�K��Z/�:��F;�jf'za��&\Y���P�����vL���9G�� r�S��Ҿ�6}�:�<�Q�1g�c�|������2�ǖ�|yAt������$r>�B��>e�^�^%U֒d}���vʀ���;"p�><�Y�
�x��3��>�m�c�b��/ ǫ��1)��?���q�kX|}|s����� �r&�]1�@'}��0�۝{�a�ՙ�����)�
�pĝ���������C�T/큅}2Um�}F�\BH��RL�l�,���]�,�s&�Ep�mjOwDqV��o�醄P���V^`��&� ?7��9�1���0l�S�W�qb�a��f	.��0�)k�2�W���s3J�EB�[
�6I�DD�l�h�T` ���H2,�����+��d<�����G����:-��v�ؠ�w�]�?8�]f����8��Gm�����@�s$Q�����/���(�_��^��۬�
��L�dc_2lb�ya 
G򖵶N+��
xV�Û�8��]�E�ޅv;f�g4͐ �Ůj|��$���;j�6���4@瀯�G`��(>8�;$]{"�̋s�`��tF{.|���פ�ԡ�ʳ�s�4����+��ƪ�Y��n22��!Up�?���G���-�a\��$��0A�Ņ���l�Y�Xa�������)���,�*���v�2������֖�I�^d���ܬ���>
9�+�I0Q-8��b-�������؋���$]��Y�c3�+0�| 0�̾����.����af|�����3d�����G�cX�����aOHƉ��O��St�>�	`��QK�z�����bEz!C�aE�\N��a6$|����T%���$���6<���6UxAA���ß��~��1�d`@���6��C��m�xwz�u�N�9J|����" �<�{2��=��̼ ��Iu|�q�⋥����)�2�^���ԓ�Ù�۞��W8��I�И���Ac��t^��9�/ �꘡M��=X��G Ƃ!��E�H�Ea�v���dԦQ�u
���͕���eV��jy�D*�6J/$����NX�9�Dq~hc��´6|Հ%���8���6��B����N�:RfG�°��W�/�����Ñ�a�=�!�Í��r�`o���>:�$��c��F�A�"�f5��H[r���/����QA�k�l+ ?�����d� e$�wU
g�{t��D���6[�P���~�\��E֞X�[ u��ga4w�*%���5Q�`�0�3}���a���j��R�����"�� ����_�z^g��F;�P �mj�H�c�W&�kT?x��C�/S�l����UH������n#�m;	,e��}l:�hZ*��l�����TobY��������"Sًˣ5��㊂��ܺ����E�[��wY4g�f���B6�,�Dj�wz)T<)c��4�UlEv�,~{ö�\�5�U��O���z��{��<K&��_��t�e����
��G��@���sHu�WSE:�q���gc�:�u'�],��9v;��UZ}�^.d�$��S���Wk�������ʔz;��I��2�r���jfݫ99#��GuZ��)�c��ܷ���:�8�pI��Y��~��:���MPc�٪_���XW!�y�Y̻gEw#�"ɞM\���)��"A�A24�v���ojܣC2�/L����N���܄��}�z3!Z]b�ga��tw����s�~/�" J/5���l��s���/�ʹ��㧾�=`a#��g�^�H!.q�u#ޢ���Ց��oP��8N��!�J�)��T�p�O���s-d�:Co�ѷ;zͣl��q��{]�1g���ϔg��<, ���-؋.��P���z��
�o-��P˧K��p��5��G}Y��{ƈ�{�i`�^(��TM�]�aPj�05�|s7f'�m�|��Ǒ��"�!��AM�l}�.f�9�O��[�Zv����`0�������Z�-�� ̡}�Fe}[J�#�ŷD���� ��59�A���y�(�ρ�d�u|�!Hmݦ  >͞F`���$�-�>nmW�g�j3����UNְh�jL�Ծ���X�M�J�eѴ��_)H8$|�m6��!�T��Bw�Ih�W=���Η�N����Y �A8�v�}Tѫ1anc��C�{u�_��?�G|E#�45�P�%g�r7t�l&�;������b�����I^��1���^BII3�E����z�-Zm�j�W1������R<j�׏���l��"�to�0�l�iK�����I�k�X�7Sc�3vpu���B��±ˊ��VG=%|T `���h�Vf�z��i���<l�!�<��
\��(�j�v� .���&I���!������U?&"���T�]��GEEVr PV��C����}���)D�[*z#=�U:?����J��4��F�]j'��/wI~c�h��Ë��bf`��"b��cFrv�ﰡ��J�չ�{+�B� (����|�����/$G�h�ͅ�/ѝ��l�CPݖh�Ffj��1�vqł����@��4�@�F����%������h��g�|큱�F}%L�ؗ��;�l[SG֟�o�Ĭ��d3hL?�?�?u�������ؓ�|*� m�/���&d�M�km\7@ʣE�_Scwshg�5)���O:[�n�۫}��y��]rב�a0�dʶ�4���m>���) �G8[�p� ��V1M�5�fk�wI`�\�^��]�}S�qW)��αv��p�Z5ǲ�F
7�l0(7Ũ5�u`y��9�iB��W�;��Ҧ:ߤ&�
Dz���3��ڃ/��T2�3ie��c�b'�rf,�l1 ֬���lħ�X� D����͆�s�^h�2~t��vE����1��_����񮱗�d�3��R���\/��"#��)�1�
��>��O4?�a�\ 
����]5f��
σƌ�v$`O���������!.,1��1!hV��$w'��C�(�{�$xE+�8��ø8�c)z���VH����5�E�q̔-��0�U�x:(w~d�eQ(��Y��V��l� �D���7����^�iz�i|)0����U��꛿g���wV~p#T�y�[�2�!i�%��Ze̠�ܶ�MB���B�0�V�~5�@�{�'ɋ��z�y����svI����7�E�O
a���E�F:#D!��8�Lc�ռ�)�W�*.�߰x�I|?Z*�Vb{���}V��U>��1���4,+��OQ}5�z�����ӢA�!:U���_�
|G��feߤ�+\�p��G�$O�O� �0��=� �����KU,�V���L�/H��s�C6��FA��[�礽���wA~#׈;��l�/�Ҫ�i,����U�C�?�v�r��"X��(~���9p}�e@�U%PvTL��iW�q�T!B�poyx?����F������wp��ĩ�t�t�ղ�[��7�v;w�@OI(�J6k6>���O��s�ZW�7<������-�i�`p��{'�s� �&�]e~���A��`���|K��[���tL(�-Y����w�8
�2"_N ���9�e��{)V}��9M�C$���a�Z��Ⰳzxj����ފ�~=5�j�&�=`��j�ή uX}�Y�`JA2;;�5�ԛ�ҙL����7�<2L��o������f&���ҙq�D�<49�1�+E�;
��qt���h�#s+;~k����'�2�j����O���v. -iC��E�Y"�Ï޼; a�z��z`��aq��b�FL��D�3(6&�0 �KF(�`b����}g��|0�w����P-�L�&=~+B��>��X�ċZ���H��%��o���mܻ#�E�74?�Y�M�������c��N����.3�t�rc�O_cC�rv?=����^���>�m*�� Z��=V�]iA �LwOڱ�_���V�3ڈ`0��K�_��Zx� �����w���(���ـ��@v��	^�rN�R��b=d�%�sӲ�}:�l�}I�#y_��Už>��ŋ���G+���Ķ)��K�(f8ɷ�N��h�>��L ��:�~�=[8T�;�_���h�*,˰C l��X���)^�Ȱ���G�ғ�8J�@�L�K�~r��]S��
:����T�F�u�|9�}�2E��+e5�K�\��M�����	�|�'��Bo%�E�}l���dG�!ޗ%У�l��ii H��eǫ-��%���l�_���.�E�8�u��>ǨZ���-��uM��2
����Dc��]�YȠˤC�u�_��4�hi�=7������Di"�-�Tby��}�̀�F�M� �Q���7i$
c�N��&i�r��RTw�,�
n���Ǧ����ˇ��U*�ּ�����`�J}��a�ɋ����A	ڀ�����{B��)h��̎,�v,���8.��x��Mr�'�N��
T��R�*�	��ٝ�`|��oc��R��x>qѲ���V!l��<���������nݞ�Yt���Ğ7}6E�D�}��e܎���[�^c#����a�FP��CFg-cH�g��V;�4��H�j 3��-H�Ų��PdiЌcY�����L�I54/jx��;�׷\��~��][�J���$AX6�`�6Q�#��	��~��t��Ls�t�1��V˶ٲ�RĔH2[�u��=�jҋX�w1iIO��� �ɗ����R���U��Rn���6��^��8\_�����Bz����9M���a�L��]��H`��y�s>3,B�.��+��\kۜ`WW7�� '�gD��2��6��BG!鿻vғ�эR#t?�q�,�PB�mǕXA��I�I�T�p,	��y�i�e[��}%{-̙>A�h|UF�����N�� 쑨×����Q��ˇ��n�5�� ,�ek��̰j �%�t�i�c�u7�(/� �{�f_�_`� p[�~���|�K��+��!Xt?��y
U������e�[�����;%!"�\�!�8�ק����E��ߗ�u���KQ��@��6�_.'�hف�z%��{��C��B��P\*y�}��=\&4nz�\�o�a~�ui���K9����I�[5%�G�]�Z�Et���T� ]��x�mۈT��\�Z�bo��C�Xi[��Wv'����'RW��W�%^�hâ�j�S�㋨@0��mL5�c��	�f��w��DC�Ota5.�0��h�(��+o��Ƌ�5_.�AՍ��yO��3j��Ke�:�C���]�X%�&w��>��eĺi��z�C��ej��9_��C����D����>�����uU�@J<��";�@|>�;Ā������1��#ǁNLW����`A"�IrpQ�KێU_���١�����(sS�����N�RU���l�Ί�bw�m{�7���i�dLX����-���=ht�E�����=��X+�<2�o���\�T�������=�7�6^�
Y^q�K{,��8f�H��n����<�zۿ�0�gM��	�_&��2Gs�F��/\8�R�D���A��i��<*�^�rBcSH1�Lz��?{�c	C��ǣ�-S�7iF���<Zҡg����v��#ص�SD�k�q��;�,�pc�SD����lnz�89�\�h�=�Q��p��t�R+�)C�Y;�U���%�����%~��2Y�s(�Q��E �0���ي�_!|��c
J�"-\�B�
�?���%�G�cm�%��3�hr~�x�9ż {��1a`�t�/�[V�Qn������T��|z�)��9�q�F_�O�]zf~w�9R�C^#.��(�>j��o����qr��	���5D���W����5��~ӖV1�ݔ��4�R�h�G$U��v�~/űӻ�Px�@=s���k��&Ϩt�/y����@��a�X���B{#��C���P���n9Or�$���o)#��Z���`���5PVV�����Qf�xi��m�x�q9m7�uf�,�5�`3���;̅�8�>��!>5�&����Z��a���>]��@r&)5���w����������)O�n��tL�U%���	{uş�}�
�1�Y���$��̀��A���b���:*�+Q8�A�{$��#U)]�]"����7���3��'�=x�1�M�D����G,>��-J��=c����N��S����y����;�S�_Cܡp*͒�+4��_``�!X�9Ț�h���[��2c��M��^4#E�ߗ�����<~��� ��'��M<ܙ3��Z����n����M��R���쥏�.H�H��[�����Y�(��؎�վa2�L�q%]j��)��7�jQ �n�pG�c���'ԫ�`���8-^I�/9��Ո�@k���U[A}&_��~Q�d`��Ɓ�R�`�I�f
��j�)܎4r��@��LP�?:g��DN!e��o��ZЯʫ@�{H�Upʯ��YQۦwڍ���!1�I+��@�9�DR$��	<�*�u�7��%�	<$w7�&t���q~���X����v�@�c� ��[�W�v�lQ�sҀh��<!}֋��2}�S-��=�3,�9*9�X�3��~,���(�$h/��k���K}�Gr&�V)r)��UϢ�H��;�,���J�j���jQj���ġ�6�T��Q7{���vF!�<�qy0/B�K�6ē ����������;T�MyV�dk��5k�;hG���9�
#����w�	\N>1��b,ؠ~#9����t�#H�1>�Z׊��O>��ߤ�.�����r���I@��w���b��������MA�ŀk|k��ݭ ��7Z��O(]��+�E�["]�Sࢭ�|d�ζb�5��l���"��A����|a�,s�W��B�D�ۃ�����0�N�p�2�xC�s}?�T�0� ֱx�s�L���[��f��q��)�q0���V�l�v�����l�n��~q���c�Yηɲ�Cz/��=���#Ӊݻmt{�>I�帝%�#�"q�SiU�Yj|X��<���[H^3ֱ����>$�<��J��k�Cj�������,����D��F���D�O����-q�J���}5��P�SZ��8!�W9�;9��8�z�����BV����Ͷ&s����2�5]	Wt�w�/��&qD�^a<�Kuөk�D�&���H-�4�X�ݏ���x���Ρ�x_g�r�&s��^I}�!NaX��x�a�<�����Ʀ�A���H�P	G����� ��Z�[	$�O�j�4�i����n�1r����"�D2��,(l��r��슟����Q�:b�����H��!|��Ď

�t&���(Jq�
 Id6y�~��$�:��_��\�6��
�VY156l����\��J�t���Q$�Z�`� �1��D�Gw:��d�bl �)�Ɖ@��;I?ٶFWq����ܰA3���9)�D����q�9B'���<^'���~t[%�yl�*ݙ�:�4�,�]{F�0�AyN�ǘ���gaLSD`���-s
����NE}���R�e�����d~�k����C3n'��]�����k!�U����[����3ך��!�L@��5���8�µ���\�W`�~!�=�C�Q	�#,#H�T�o�<K����]6�� E%,	z�x/O��D��'�+���)��}<C��lneK1�ꀴŅ��4E��z�lU1ߑ��!$����U������)��ȍGAN�7 �]<qh8@�.��u�[ͳ��I���� ��'[��'�Ǒ��>��N����Ң�(�J����+f�T��F�T��"��1�}�_�{/}�}� m���>mw�R*�4��X=g��S���X���R�CUtu̬F̮D��/hwU�2C[���0���x�ʽ~
$ ��
��>��Y�����y�#7k��.����6�Đ2T��{��/??��4{ch�+���S��	�1�-%����.��{�WJ1�18�4�i9�F[��I?=p+n�[��4`�ތ��]JAo��yfl3p�q��'�FiX4>�)3�S�ε1lU����'G^��xM�4�`{Mi���X�㚿辻�h� �8AZ8b���E�������c����W��!�q�O��N����Q�P>�'>�܈�:L��lR.���P��	(�j �O:}�B�(N�<���yM����-��^����s��B@Ђ�W��xS��Ձ������ (B�/�ȟ7�C�(<�
����},�����O�x2���T��B
� 60�Q����ڱ�t�,��xj3G�	��q��5��M4����N��Z�������H�5W�y�*K`p�%#ڪz��j7���1�3H1�d����:�w�b"�U^��'��gv�� �lwnM�$J����@d�FJ��9�}�C}�S�@��>����r7,���_p�䰠��*%�>���������:a�*�llm�R�`C��`����db�@�
��@x�pEj ��9rK#W߲ӹv�b?V��؏��)�T�����1��q�ћmp����F��|���%Ģp��+?���fy�eY�e��`;i��������Q�"�����y���4�xD�e6hy6�vN�|��p�g�m��[�WWQ)�{�vrvH� I�-aA�j?A�G���}����@���X1����'v�^��BsR�F��4�?"q�����I{(�)�V�cDe~�mPV3m3���]��;�Q�!�<8DՍ�Y)��W�!hE��)�xd��]D1.� �*ơ����hn�<�I��8�,�R_�YMNJ�Z(�o-��
�掛)�*%��$Z��MqD4�6�:�J���=s{�$���G����og�Qġ�N����迍�jj�e��:�qt,x�p�BD�� �>�̙�UR�,"jB D�$�E���r�5���X��1�e�M-����}n��M�'�N���\j4�7aM�)hZ1��sԚ6���:��C-�y,�q�E�D�Ӎ�5�u�y�����Z��I��Y�J�!V^�)�B�M��']ĕUp�c�x�p�Ś�-��:�VP�G�q7M�{�`I����`x`�<�=�v�v?$'���y�t�h¡ďl����oz�U�K�^b!��>�7��= ő)�*sq;3Z�M@{Ѝ�u�m(��
�t�[&\(�y�z���ն�N�2��2�Ɍ�@���t|��X�nӿG)�����ȿp�D#�Qҷ�� 2�)����;v�@�.ѵ�/bɻ��$\��3��'��U/8���2Td���R]�Y�%��	
�]\nS0��Z��XG%�q����T ���R$%n�i�7Ж�L���rx�+W;��34;���3ܜϊH#�6k����ʆ�/�L�������+�
�=ˇRh�/��V5��av+봓��la%���˅w�Ġ��}.t\��a�d�o{z��V�@1W}_���~i��e���9��V��4f��kPA��^�aX}��p劋̑�^��k��3�JͭT�mS���~�j��+%V�?A�����G2�&+�/������k�A�82`�9Z�ihDՑRn�ެv�b����p�^?D�"�����6@��$\HX�Q�d���g3����� ��b<�C�	i�_Ķ�kR=~�:[�
����e�uT�OJ�в5͟��Y\�t��K�R�;2�X�N=�z���)"���,X;]q�(�w���;�B�?pd�Bct�:2x�B�,3wp��f0k%Ť�ZQ�� {�V��>�"���|�&�4���}Zgf^��K�5-h]�m*~���k.$�����{�6���&%�4�G�Z�{(�e�ZM0n�q\5/��BO�+��:��ݻ���B����t����(#�o���_���;3��C�3$��B^V-����<��A��(�E=p���/�c7F�nrS�z�����Jv�p �C����M�B`����|Ϣ�5E_��[�r��Xiϓ����N�>h�X12�O�,�{��uճ��EAeP���cmi%�Z��<�C��^�
"鶗�����k�S>�����cL�Ǵ���aS���`��{8�=`�\-�F���o;�����U�
�d�8(����q�"�fQ�-eF�c�џ��%�����?�A�-X����[pq�bCq9��bV�\�@�i1L52/9+_�0E%XccoډB��ϩ"e�衰�2O����x�T������
\�P��Gp1���*����PX,0����HE!U��, ��'W�$Sl�q�>��	�xd��ŏ$](�|�*��:�*CM�g��V��*y4\x�^ʞX�J�^ڈ�כ{a�^wb�i�]��+:+_��j�nm��/}*~y�,TQ��R�\!�(sl�Im�^�Ƨ��Ԡ,��e_���ͥ���C ]a\���'��۵�4��#�d����w�,�U�8"'-�Dlf���l��-��&|��i��HS�����"Z�%����4x $x�5aJW-�I�Ж)/\�>��#c��>����ZE�i�)�hDf��JZ<F�X�|���ң�+�W�bX�7��lԾ��5��#r��&�ST����>:f�.v���&k.��*e�,�tK����^�����N}/4T�ҙ��I h��$��d����EI����μ�m����=��>0x:>�|���G����oY 49[j�|�eq����H��z;������?�+�7d�/N��FjD"�]�ǎMC���1��G�A��[�vX� |';�g�з7�����h���j��_��p�g�p-PM7D�e��J���mn�T�a����9�kJ�}��z�XW�$�nEԴ��!]��C��} iK��$R� GO� ����[e�W����Sw�%��em�];�8U�r��c�3�qg��Nٺ%>�0$:����b�aC������� :B6`����A����pCcn�E�LD���k�/y��bؔbQ����}Wҿ)����ܪtI�ȣ���]���Jnv�)�]���C����66<�]��4Q ����%�/�F3*6�n��]�*�)ͳ"�1����5+=�j���_��l�����4�}��J�Ѻ���5���������K�Q�쫝�o�F�Tz*�w�ڔ�iI���dA���WzW�}�G��Nk�C|����|Fe-u��1�2�$m0q�i��k�2�,��3hL�9�u�g��ȿM#p8�:NV��H�T��WK���J�:������_~�,��^��9D.�+��nݰ�r�XsnG�@Ω^�X��<���VJ�}�	��wf�D�eo�^yL��9[U%�6��j%=�e���,��O	���=��$�d�{�`�Tk�М�Kw ^u:�n�����Ĺ ���'t(�wܺX1�4��y8�5����@������z"�����*��M� �,¥�P.@�ۼx��͗(������[!3:W���[�1���k�g��3�^�ǽ�ɸs�sT�9)�aP04ׁ{5���R�A'i��J�.;����]	n���%��~�|[��{R[x�̥�O��?E8��D��+��VY2��k�l��`_�~>^�M��i|�D�5+��p.��Q��!ܻ��*H"�~o�ޮ����}�έq����2(�
����a4b�=I\e9_d���Q�`[����_����ԅ)��Z���� ��`ao���m3�_�zh�TɌC��xC@�$3\�6%"9��Yn7F��׏3e�*����o���t�+��oFi����&c�
�P�ۡ���=7���`���g;Nv� 6��"��zJ���n���Ӧ4���e���e��"/�Gd�w8���	@ZԧY,\L+̑��A��[�S�Մ�ٟK"�aK����څ��{�^ɪDWv��>"���)^Q��H��#=uYY��]at��+g���8"sD~m�"Z"��L�K��kN�i��̕vJ�&���=&�$ s��O�G�u(LĠ&(�����x��x|ˬ��� �Ԍ=-��z!�v�r�B�-9�߲xA�J����ҿUl�O���
���?��c�8�Z�m*ȸ#}.!!�{L���z��_g[���~:/��[x���v7��<E�f�S�f=���]���Z������;p������Br���^_m?��C����cX{���:`%@�1��>�Q��PA�� �^�@+���a/*>^�\��Z3ߺ����1�`m2J�y��(]YWC5`2�n^i'��{ێѪ����vI]DȰ�E�"��A�p�p�f,��j�֗���J2~�L:)����Rr��v��+x�0�3�(�Kh�)�Zݼb�cЭ�4Ӑ�+�RX��ޮ
	X��Mٌ�a�$�{!�A@4uW0��k�vitS����)�n�J��Ͷ �Qq��?�m�t���D���v�B>m�Y�m0�"-�mMV1�gX�w[�^�ΡnN��,Qq#�e�T�
�b���^�苆ұ[~r�Z��zX$��M���"�.�&W�،����������QQ)�.�|J!f�?�
v�G� nS\�	r�)�xI�]\{���ʞI��S<ŉ7��1���帝�[���ҽ�F�����Q�PU���e�y�#�r���&Q4����b�uX�ѫ
� LEIP�d�?���2���U�a��`6��xC8�q��]V���|��!��r��YZX�q��3A,��YA/^� �SF�8Cڋ�IGB��ז�ʥ�����7f�k�1Sr�maxq�f֊#*�^�ys|y�&� � ��8��g�54KG�SE�r�� ha���Z��8ᫀ�-f;]fe�m]�~�O5_��H,u��|~���ؘ�2�E�C_�R.�	T�k�Qۆ�e5��D	��j
�Ѝ�����/x�yV4'}�����6f����\�m5�V\F�6�+K�o�['�wIT�L0�b�aG�8�J��$5%�*==X!*�Đ�������j�<!�d�50��=ǘ�o��*�b_��P����>-A��x�O��b�s{�~�P�D�Ak)]�U��D�(	t����Vb�x�rT6�4XɏD�,W����o���5�Py�)�	�������j��&�֒b=�����͓������)��r6y�q6}���t}>�k�I�<�bQ�
��������^A� ��CH�ZO;���H���W��͘�7�O��W�����(�TęR����Ne��D���]	̐s�ɵ.E'��NR2�o���,t�,ZY�@�"V%]ݴuΘ�B��MZ1�U�-��A�T.$����0-pdMh!��< Q�(a�hstr�
1�#"�ڳUpU������u�]EI-�����\�%fM���rٗ���f�Y%%I��J�����d���/S���<��*a�EV�O�La5��������rO�@�����;(=�<���ֿ�u��J���r�ךG�'�9��w��_�0��>�����6���}-N��B�qe�v��f��~[)�4ͭ��>k��%�N/��V��@7�%�Ɍ}k���5o#G����̗	)k��0���F;�k����ܠ���Xi1��?k<&�Gza���k-S%N��:�� �����Q�H���S��>���iz����^��g׍�/6H7t��!�f��P����D�-�ל�����pZ�Vc4+���E�xr��8k���,Z���y<�o(�?�������=޵�g�ئ��_9uĒ} Y ��q���f߉����S����蛴
�f�u�$�k*���O�貿�S�q�L��?X� �
4�8N	�e�_��-��z��L�����?[��	=#z�ư�'�HI/����������|��#;ڻ����1����͓ޖ�@��U��*�y�Fqĩ���H��E��B����~>��C�����p�{�-8���}=5������_ݼm�JON�M/&~�i������b(�p�]~��ַ�d*�M%��W3
k)�a�7�R[6��BpW^��S���)d�M��<���#��8�f����j�+y>Z�;�V%-)_�7Ht�K���%�)1?�E����2�?��k��~>��.=�=ȳ����-^����B!��s����D����ml�G4����{���oI�|
ڰ�O�ql��R(l�meU�(�Z��K���{/@ޥ;:�,�s���~�W���W��(t}��,��9T���J�l�Ww��L��9%Ue��K�J*Q]`�7����4W�U�}�鰀�.�[C����>}K�-�mMgU���/n#��U�j()����������~pe�+�ExrF���Q����NO�G�Q��EoJ(�`|DW�R<_�1Lk'��_�q'Ɂ~5ƌ+��Z�k6�8c� B�+a�8������ȧm>S�9YzA4����K�+M��)�w��*�&G-Ū��"��\3s�N�Q���M�l��g&��� svk@j�٣�*��UUV�/X��pԢ	uuI�l�i�Fq0|���o=^L�e�_v�^���`�����VS�vHp9ZiL�K� p��Hom��79��Q-��+�v,��Z1�e��JZ+�k�q�����QVE��s�v:K��������j�.�&���f(�JZr��x\����*Ȁ("ʈ��

1h���|�Z�M2�X���C{��X&����X8�tT�TK���v�c�b 
ſ������ȿj�����c��ut��e_�o���=��6��7��XWЕ�VT$摃��A�NE]"+,ݹ��>֩Zɯ�V��x��)�_cm�I<���6��e�_��=��wA�@������>(�m|��*����P�P�䆟�dA`f&1��Q!�N������N!���f�:�J�´#L�M�	���v�ۍlc�*	��̈����j�
\KW�7�L	]���4k����8����m���-G"z���x,	{� ��͠�n�
t^|���@ -�ʯ��C�s�`��::~� ��]��L����p���_I��sl��!֡2:K0�?
��K�e��w��_h�u�Zzz��G��	$݂�e�dvᦰ
�J���8��7����A�4��\"N��8T�f�u�W�
 ±^�z�kw݂�e�(_Q�F�<���w\�00���;�z'cC�u	���&\�P=Y����>5W����ܱU�׀CQ/��%=�����/Xm^�`~����y(̻4�Z������0�^��|[��j.�N��a��/e���_�M{q�C����ϕ\�ܣ}r6�+?����.j�0@ :+΂����������g�MZ�Q�&
N�7�33�S�xA�9�c�)�P	��}WK�����hhp��C�Ռ�i�]�9�k�|ܻy�LS��a���B�Lu6��(h�ڼ��q+uq����ǋR�	J`bǄ��Ϸ��1�h9I����4]mĠuy�SA�0��2w~o��i�S'�/`��|�@���7R���к����JD���ihО/A�)�ڱ�~�v��}�6��ڃQf��E�(�x�6����;Rb���'/����:�#rA�8�wg!�6��#-f}d\���A�:P�x�݈�C�<=��&hY���'d����c�����p��U�UrJ�wp�6J u��H�`i?�©{��W&�DO`Ֆ�	�'�3/ᅱ]����b�WCT���;C��*��LNڋd�9<�fBc.Rj���2U�.�ȼ7ǎj���Q��?+�Ӫ�A�t'i���sTg�X�$��I�odNrL���L1��8��+��9Լ�'��� �n�7��yo����U�ж�/��#�J�ݎ�^����c��q�&�z٠�/�(�s�w�([�JWy��z>�u�U㤷E � �Q��[_�� S���*�������|�j�����[���U�qO�VX�t3�:��h]�B�je�؝��GI:��=���;���,�v{��zf��#Ÿ��1��H�0h	SP%�%�]71\��:i�$y-�g����� �������?�j�\3r.��l�F��_�jw6f�����?}h shs8��,�,7�<��D!�k��=~��,1|��w��������T9n��v�xi�p�D��!���;��������4}����W$�r��2.����F��+J�g��=?��z�L��R��#�=;y_ws^�H~�{���[�3%Tq�~%q��֌�4�zV~��L���	2��m��1'+��|K6}Xi��К	���@?���oq�چ�B@'ˌ�G��̹����_S����6�"��#�m�����<B�	���M+��1���V!A�ϥ��s��nH�YMJxz}�sv�P �>_�ʦ�i��m��0�y�e�_+jպ����L
��!���>m��׽�&(�Zc�u�����A(֠d������FǬ���f�_A����t��e�wa��T�7���<&�N��6@"�N[F楕�FY�b�û��'C)#	�Q���(�J�'k8��b�|D�Y�<��`m��/�y��K���P/~!��z@)�l��Or���S=W�<��h��Q�L��ø�����~�b�a���9�������^��z��!��\J~_>�,ײ7RQ�1R�7?4xĨ.r�D�0�3!��G1�%�ӝ<��J�1�Ez�&Ra��>��Qv�*?��':o�G���Cx����aUuC�x��DJ�ɳ�m��b���(T����7yP�M�U���7.��"�HK�C��\��Q�/�^a��F��j��9�-�i	�f���I얋�IN}e��i��`�*���ەW$�P�Z�D��Yت�m�3����ǟ�	@�t�:��3���.�g�XGu8�s`��b�(�!h���D���873C4�A�u�:��I�$�ǃ� &�@�Y����M@�3JƎI���r��h�Q���9=Q(z�߷��׿A/�B��T�:O��%��r�j;����wWw
46,HK����UPI��I~ ���eJ���[���4��|
�'��"綷�f_�4}�5�%��E.�o�D~���a�nQ�|y��Lts[����[�8:���9�e�3��6��a����SE^�>�Y�Og�.��\���5 ������鳧�c�W��aq�C��d�O�B����L�N��v����rҾ7;�W�(�b�<K���_��DW��Jh��$f�drZ�	�����f��<��#Ȍ��_�Y�B�ߪ0�օ�-:�=y���7���U8�&dOj�g�����6"\0(%C�U)���*�h�<�o��V{�h�6�N������l��W�󪔨�F̗��sAa�K�S�����1S�|E�f�@3�Jx��	��-t��,x�:9��P܄⋗K�~貽c���h<�&�@3;YByqn�V��߿-}r�EU���T�w�bY��5v��%c�iz�NP=��4!����"��5�c���Un���:
�l��&LY�5�Z�58 P��������jԸ�2����oj� D���~�od���A�����I��#��L2��G�O��f A� �  S`£����]0\ؖ��%J8,�	  ��m��0�N���>�= �+r*��S��7LlŬ%t��4b��S��%Ț�� �?kۮ82�9eZ�Tn�" vj��j62u��PHȯ��xXވ"�1��u��4����� �'U�����{��9�.���}��9b!+_..\�4W��8������@>?8 \}�\d^!��5�F�33�*���Z����PvO��;s��5u ��M��ɌY�,�/�@��AQg�:2�,?�L%٨��}j�R��.���3|����E���o	 T�\��D'H��Z�V�:���yxG/u�	#Puk=��3��{��,.�$�-d���R����ic Z��l��a��z��d5�G�q����G^mv2;�O Z�V��<#&J�i���_
:�i��>S���O����qێF��=��s�G\���"�kDmL��&Ó�@���_��/���e�EZW�1,�q3#����c�
ǌ����^gSa��Y���h��Z?�SH�'�C-B�DW�_G���p=o,�0�%��8Qa��؈�
)�t��צm>˒��v��������+�HՃ��t�%��[@��i����wMe���i�_���-����:�/�x���5w��HV 6�����]3���z�v��½�"q�F��A���Xo>��Y�(���t��d=^�"�0+����K���;�IH�D����	��l�߹�S�]\�^�\N��a3°]�c�x"���&�ZrL��#X�Śu1T�و�#�ZC���>bT�aHH���V���� Sϫ�x*.S@��^&�ֹY��Q��r�U�;07�u#UŊͳA��$[©Ĺ��ƍD�2'��L�xp	yy�*��e1�g�=f��=�!��*��]��_/_f<�wd-�	8u�e�`�z���4��D�@��%����7��s�#�/`�_�X�9y��Ͷ�/~����{�U��gY�_��h��2H�U��q�����5R�5��]ç�� 
!|L����[�:���`�9cҒ���i�S#0�4(�X�$Ϋ�̖�)x��r�a�{�X���݅���Z����T=4H����&�Bb,ץ����3ah�g&����Ƽx%L$����zz�B�-�5�J)
���� ���;>��nxm���m�@�Z-�Z��(@i�(&�PXt���D�ϋ��xO��g��n�1S:�~�l�@%�X��U�T��44�CW1e^�eA��NV���dR��K]�5B(�'r�)�pw̵[�]L���Sx�y,4w��L���׽&�5�	��E�J��K����O���.�ܰ�+q]�a�ɀ��%y��k�c��%��s��U��>*�!3c�/������e��Jx�uu��$���،��|���׵ggO�M�^6?��ݹJ�rSܾi�=aj\Wy�-]W����,�Wh�����JY�{T���ڄqu��G�E[���/���A��X���JA��� j'�b�R�z3�%�w��vH�E	v��#�3;z��t�Fn��-bR#�sfƲ[2��p$�X� K8�\�fy"���S?ͭ8�]�9�D�(A�K��H3���������y�*��Po�+6�Aj�����D��J�uưsޖV�?�l6���跫��f��'%pi]�-U8<�~ȇx�k�}���6�������>�_��HY�� q�-H����Q��C�6�jƁ{�K�~��� ӂz&ȵa٦�03UW6�%h����q��*%=١G����	�k'�^��hN�x�Fd΁ܺZ��:�����21�dKtw}�II�����w�d��h�Ƽ+��� [c���BDWt?�@�.w�^������M����끜��lP1�X{j�/ɨ��^�ȳ�"/}vHOC�r&�<+H���l���9����w���1~ǯ��8f"���,Y��Mvq�v�G��H�!�����x֋E�p�%P���-��lc�#�v=lQ��L��.�V�C5D.�@���j�.;�P����!���c�ZV��`�5�ѽe͗a;ث
*~�RCݳ!.M0��si�y:�d����|2�.�D�?�ןnI���X,�*2�H
����Y]v\��C�~m��ū_��|L4��-  p��ATX97*�h���K&8�@��~*�O����X��L��È�|B|BOYbE*)%6��lu؄�&!����D�h�%B��~°�nV��������v��9�E��֥�`Ap��bIX?�ҭ3�Q��d_p;��ۍ����g~SV�&��IIn�2tc��i�t�K����`���>=��5ހ��В�}
9ͅ1�l��Ő+@��tg�G�]؛M�S˾���%����_�~�w�o'���X9���h�qs�� �W�ޙ5���NɓzW�
�i���Oԟ1�7�ʺ��F�';
{��'����=@���Q\|����Ĕ��)�Z<������}N~�[uP�+��u�pMpT��?����CS��f@.��a���'N^`��6	�ܪ�����0'�j�fA����SF��٦.G�/�͔�֛�c�c�bIn��Б��5��yuIYߪ�
��s;��xc�t���nM#���=����j�	����lL�G��z����nf���3K�Zd�M:�ٟ�^�Z�zM&#���<O�w�t,���u��w���h0{X�'�N���k�\��M{ҧ�[�5�M�gN���A,���NR��T���+hk��K3?63&�P�?2j��W�gky����	Sw>��̍��Ai�H�1��G�y^&�[C��[���T%�YlfC�"%��Ek�b8i��p7�!�i�G)�k?��:�u��2m�0�Hi�k�bS�6�Qi^ ����M�,�UOc ��9�dB:��~��G���8A�5��pS�?�_6C`��.r����S���y��pef{┭�l[�VД+���:H�i� �Ⱦ�������0�n_��9U�Մ���:���S�\1�W<��d��	^5�t5��Yñ�Z�"&�!�yݤ��q�&�c%����l!"4��t�V^�l9'�ZF��(���Ø�'BM�y0��;q���<�Cr$�L�Oo�\�{��
3��G�0��r(.Y���R٬�3��E�3MT<	�����iv���Oè�c���U�ɭ�Ah�ՁD�A�^���&��0������_헌Jgm ,���Ҩ�/�esd���(�zqA5;��7���>��� ��ވr��Q���C�������p��G|&wǓy��*�&��͘�+�k����m/'$�r��
�%�oz�)�s	R��?�A(��t*�K<�W�� ڡvڛ��P�N����33aƯP̼Vä���.E�Dc�ƀ�=�j�۾8q�������܎��<rt��m�O0xs�(�(��.ڛ�Y����a�+���(+�l�:�j���S��idp������o��ʭ��$�H0wq@���'q�R(� �9�T�'J7z��N�4�v����E�ނ��Ak;.5�VGP��u�����
�C��!�Fi��U��;?��U��f2&pIG1Iƈ̇W3|vG=�*(��'�E���RA��$�{a�
��A �ɴ�Y�L�M�C�~����� ��J"*9PC��ᡔ	GL!�!��`�r,������rs O�ʎ�`�a"�����[�-��!�OW��\mK4)���jRaN�W: 8[B�MWiS,F-�I8�4o����
z�`R�����3j �*�ߚ6_�\���{�w���7z��웸wKX^���Q���s�.�����=�g��w�/���M�<��4�w��K��y���kx'�f��;<�-�ػ2�Aa���O�cz�Y�~!~�����1�E�mL�R�n�0�U�=�g�]�q$�袑�3)TQE��������� Ou���<W�1G���A�rW��.�XBSLv ��S -˱��l6 'ǇG��� ��Frhp|J��3��� ��i�ӣx�9s
*��º%x�ͪ��{ZKE	���ؕJi�U�О�ЇFL��V[��[��YI7���}��L��CL�C�i$G�;!fb�Rr�;�²���W�3�6�=dnF�]�-Zk{CAjC��E ��Mb���4�(�a�/̗囧E) ��ͤ��#pB<�~1�����э<�<�|�\�8�Æ�\�߿�!0�n�L��
iջ H�ďC��z����<^�$����<�A�?�\�������]�X;׏rZ
�>CmbȺ2�n�y4�Z"Z��ɩ���U�HM7�I����HM��~�t��Zk7�
gMϴ�6��f������?�my�j6ש�"~��}�mUTh�b =�{���t�(�꾻F�g:L�?!���dX� ����	�ڷ~�Ɇ���7F�.y�a�D�>��I	��<��<��B6� m��$��J�6(�r�Ŷ]z�z7�f���O�\���C&��N� [�!�q�ayBe@�a�XwQ� �?���Q�c���ڕ��t"�oS�Ue=N2;��^�k�1Y�ji�O"w�r�����8����5�>�f�i1(d�F�.R�C��_�gt��_�ѿ���*;7m*w�Mt����T��'��`H�,Kٝi������I�Nɇ��V� '\�{TY��� ��9�N	l��6-����l��)�H�j̀�(O���q�D��p�-o�WP���9z�'����m�=!B�h�����zv^���^t���7&�>(�8@�����s]"��}�G�y�]B�Tsgz���\��Ȉ/釩��!D��j�+kSj�>�o��th��m_o�rFt.�,.RQZ�q��4&F�ϒ�V�nD��j���u�0��P��5'������׉<�ܪ��h�	E[����4��4�ʰ�"��nЗ���2zshf�����[�V�0}�G3p�P��� lZa��CSS�ÖY;�5ul�7�U�����*ua,t�96�T�;\��؅�Q_�X#��[։Z�;}i�jp����^�]z��]��R��0��k�D+S\��I@�u�J��ӛ���њs���#�����]�o��P�UyЪ�lP��ۙ�y�������>[p��F�~Z�Sz�)����L(��@�(@���zk3P��)�#��)I�_�������������{���a+��~��t����}���ɒldgC��$��O�|k��s΁���M{zv��o��d�K�`���%���R����e���C�´H�?V��9z+�v�1��C&�Ch�P�V!�)������8�z7��k[���|W�=��X!��0��-�/�ȍ�E�t|x_n����0V���܁^�������W�����QdVз�I�%sV}O��YK�`�D��~��ق8J<(�P\g!̀�
?��gZyr)���@����u�'!�sA�I�7'
�����-ݟ1��@�4������Ͼ�
���ײ<��ğ�ʽF�I�?�宺����A�[�?���16ᑽ�#��Z/Q:GFr���� ��SbM�����!A�OO���u���e�UObASL���kǱ���V~ֱAļ~��=��*W%�
���A��a��u��asm��*C��mib3�52�o+����`��Y��Fh��������&̈u+�/�P�����K��n���tv|:p�cU�.�;�'e,krB���{JȄ�i�WC��ꩱK3�e�/�B�D4uj3T/�S>7��9[zr|mRV*��q��Y��!�~������qDR1�Vh\��}�F[	�1�I?� �������Wh�I%�fwK����D�_�M�V�uVڬ@gK���j��E���vD�w	ρ�n��ˉ;۽�jMށ#9ߢ��3�m�:���
o]Shu�F���~��fҼ�H��C�mg���W��`;�c��H<�G((6ޤ6\�]��B�n��E@�n�(�S-}�!�)�MeS�և��#!�@ˇ�5rT�Ӻs����f�-��5+D�%�Ti�-�zG ��h662>�˖��voAe,"7S��� �9�&��o�������^�c�.�P�r	�ax�O?�͜�g��K* #������:Š�Tv�֓&<R�/tYk㇓���9�tG�#��C� ����D7��Udw`�sm"DK~�:�i�L��C�T��{S0�O����a�M�,�K��zk�����$����pL�*c>���:�)��+�/\���x�1��e��b�z>BXd[;���.+��Hm�-/l�<ӊ�D�:u�| W��OT].>�U�,cM����}�=�nBb��֥����1{������Ƞ��q�1G�f�e����6�K�b�ޠx��-��/4<�z��
'+��W}>�9��V{��ax'a:��B�CI�k|�E������� ���B��՜��nvպ;oEjiE���������P_N�>MC�}�����s���3�S�{~�S��^�=����V*��d�����_�"7����,�>�F��������O���Jl���)��xx��>ˍ?ڝ'�E�oN��d���5h^c��"��H��7���N���Z�C������}�n~�}l!��KG����w�9�rNتŲֽR�FM��hX��b���(����٢��y�\K2=��%x�)*0�����Cx�	��#�į��f�p��:�yh�,�k�*wz�����in���:s=s���1��8ɮ_����S�m�n=tј	�����%����(��Hp��K�O6R�u7��l{ ƨ��}��b�l`7�r�����9T��M��d|�R��λ�����-�ϧ�����x�l�]�(�~B��9�Z�)0Α�f(��*��BX	j��]TrR#�NM7�u����!���.�W^��\�"��@�-����[76Ẁ�s���DD3���A/�A������y���:�O,"��<���@z����&:�3<�-D�
��V�M�;��/�M,W��s������s�lYO��='�k:Y3����AOG/�R��ʄ�c�{ol4�Q[k��Ҽ����|���B`�:�{g�����������p�%�>!�
`�{����_�ԗ����s�9���$����Fa̎2��4�5@t�f��}�"l�7	:zť��x���Ȑ�A�!�;�������;�v��RP��[�t�P�	نO���ѐ�m�go}�i���j�;�a��eƺ�Z$����>��Ɛ5�P�����&|o!`L��8ɖ�7����b�E��0�.��!����ﺱ42{"Hʪ�Ds1r0��d�S.�V�~�W�6��YЁA�Ks�n���B.@�2d���D<a�,Mq��8�_�")¼���0s�v3��?W,
�p��h�� ����N>�6>��߂�5��D*��sW/��}�7Y�vt�R�����{Ph���H}�V���|��]�|+S�,%�.Gӕ]�����Y��*�Lٴ#�O,Tw� P������h���bnr�����MY��/�f��z�.�k���$Tٹ����t4��=�ܩ��� �W�qEw����g��,z���g$�/��� �������=|�aYR�_8ڔ��7Mzʮhc)�9���1��ɑ!=#��B٥DFh��	��7Hjw>�0LI����5E�iJ���]XW��
LY�t&��Qy��=q��W����� k �2�!�����Y������Bl��Vl7�IsG�.5h�2���M�{Fa5��9*˕�`��q���/���H��3RZ�����!,E�5}g�'_��ڞ؅l��KQ�ix�GhL��'ƌ�|t\L~�6{�lQ쁶eo��m�8_E���n������6G�������$�t�ս.��o�j+�m@ ����f�.�t/jR�(�`<�w���3r��*��W�}��B�ﯮ���d̰6!�;�����L�S�5]6������(���[���$En	(�����	V���4d��y�E��#?�kSX�	,Ϥ;<G\�@���(I3R��zx�"qL���])G,K�\�
J%>Ԟt;Z�wh��ueXIP�G�s����p�[�2����q	�; ��I#�ԏ���ᗊ��l�"�F�6x�]m���H����K�HN{?rĜs:tcЏsnd;&�m�?E,�������vCǃU��M�9��o]���V��k����O;�$M�C����h���J���Z��+KG����|^�5���ʥq�֊�]5U.�M�����?�ewr���ԚZtB(�jDm�u���x�~Rt�'>��}�Z�&����a�i�Z�>�0�\��߼��)3�'^��6I:���V{�F��@gٵ���,m��4?zv ����򗼙�-�\���%��O��ee���r�x��1�D`� �6h�0�����3������y����-��v�r��D�:I"!��0"x���l��[��hl9#�������m�R��LX"�W������2��z6�� ��?��%x.4�X������b4��[�t��0��k��+}��<}���t�\+�(V��F�ۊҩF	ΰHP�>[���e=!�딫Ĵ�J4'S��g�tBu�#�����s}�րo�)�[���iҜ誾��%L�oM'���^9kľvf���dm)\�ǒr&;WPho:

�m�p/�sFe��4��;B�3R�w����}e;It�9�I��	J� R5�ӑM�&.Q_��*��m�>�d����v�Bz�^4���3X�
TF��1�� a��t�h�d�"�~�=�H�7��4?L����B�Yu��a�R����=?��M��Bq�����,,�K��k�߰�s�P�e%�%iע���X�Qu��1��%;<3���hQƵͤ�c�.T+��:�Gz�'R֗�u�����9��sܡ-���@app�-f��ծ�����@�=�J��Gn��gP�$ê�i	np�� Y%���5E�W�z���OM!���P�:�7Ҕ{��),yoo4�G�O�d�r;��ҔN��W��T��^���Q*�z��)?��T�6Φ������B9h�m�7��H�: �]F��#��!��mk̔�X}��D`;/��n�N�b���8���&���>M'�x�� Z��/��k���ard
)�[|��i��J�X�B� v[`�[�(n�͂bm'�6VgX8�u�	��|��~Q)O�ȱ/�[9'�g�:2�e�jy)Sa�n�;�BE��!;p`G��7��I��27�EW<�:I���r���y\N�բ�#��(D6���of�c�`�����2ˑ�Š��Ѷޢ"F"?�͉�)iv�G�����䤋S�d6c��*\T��d͏�]��������8�g��"�R��R�	�L�Go{���{�J�ZK����1���桰��������[�Sb�1��@K�AO�mI�@���|�wu/J�y�,��������0��%{@�����K�B�<�V�~�.s�n� �d�k��qr!W)-3C�OԽ��Ӧ��=1����t�pD�����PQ�O̰�}�Ass�pJ�ED��}��7e�\uKf4�A��#��U�Y��x�|K���	�?�HW����YV�ɶeT�z�����x�j�#8��-S�M��-$�O�&�0�@��v��z�XŹ��Dǂ&>��)`����(Ǌy�6�C�%�IPĆq�X%�0�x�V}���M��h�����`�5|T:ɺ�3�ዒ�8�fe��z4�3,�Q��i��2v[��6�嬥�:Z:L�F��ҍ�����2h��P0ڔ#7
Nn�K���/?�ºZ5HYĹ��x�}���<-��$��� ��'Īe��i:g����s3oTp�a_DM��`Fav�:�@��Ɨ��� �rI4{Ï�n�� uͼ����Im��w�3���R;^��+����|Ztܛ�/B�3�21��WOF<�~��Uk%H����@�RG���t�pN_��|�hh��Q���*ֈ�`aO�2w��ޠ`��5zՓm7TdG�J�Új�[�Xc7 �4�b��/Gd:g��$2c���4q�� bR�*��l?�REq�4�7�cI����s���_��q���WC����:��{���#��h��a�_���[ ���b���(G�i�Q	2f$MN���"-�lWg�n�|����R��~O\z�FV�iao��G~�t���I��o<���+:i@6j�w�3�Ƥ�c(�6�F�Ӊ�o��H%�1����5 �����C/��V5r:�]��`kV^���;N�J'n�g�wb���p��*��$tk�\Ʃ=2�֏b�vvm{1���D�JDX��j`64-�M���, �jd��D_,+�������^x}�oI���M�M���Ee�6�s1�.�B�񟮼E&z�N���v�4�L�C�������"��e�4��#��*��P�rta�xң(����ģ�GRq�;4��
Q�%�ԋf����Zȹ�#0?3
9��ȟ�KU~�a�Āo���0,Y v�^՛�n�e#����V���2E'~!� kW~#%���Je�A��=@�(@8�! r�!dX��O��G�S����cMP��,�o �z��xǉ�uW���F�'c��R����G��,�ˈe ���(}�meFAl�@�����r�b~GQW�
C��Z*��f��p3���	Ɲi�N<�ORDDᨱ��<��b�e'��@�t�'�V޷|MB[�Tx����|��{ ��2q)p]����<��\�A�*+u2`���Ed�qf;"Acuo��gЬ��}F�G,�4mV�=kX>uհ�Q��B�Q$-7'1Gi�����)��e ��\��ç*��-���!�E,i"J#��qj$���T�9�<�m̟,�l[�̓K�-x!{Ɍ���� 5e�o�ΰ�o�*��a�������gUt���#\'7&jF�%���̃��蓊]���\��Pq�y���lP3)W��)-�gBd��B��A��E��6�j3�Y���K��^W�+\Q�{�	[�XN�*,�B��M�e�S�ʜ��Q�#ȃ�`9-��AB�+X[�uPA��ڶ
���E��� ��m�F��o '�~D>�	�vAT���e����Y�n��O��K(aE����@������^8LG��O4~�4��v;�"�K]����/e�d�]{�Ի=��a��7-yw�gKx�<����^KP~�VwyXn���� �90�����mR>�q����hz���92x�y�ɡpu[���(��b++fk���r&��ϊ����`�c;�0�j�#E��i��k`x
����pZ��_�V��@}�O����Ի<m�9��E��QZ;�Ac��M���5��i^�����r�.5���š�|�t��]�hYj�(�0@Ici�%��0@�r���l�� ��-���R��<2D���Eu�2�~u�g�vaX$+�5������w��J=/�F��?G�h�*���2k|��G�'�z:$S/:�hh��I�%KhW����"F	�2������չ<���u�$�N�;�W\�l���4�2f�w"�#�WЭ-��w:7�(�mt��1����Lu�n{/�[�������=K��B9R���v0C�*����O���q�/��0�,H�H	�I���iŦJ����`g�P��[P��?���f=G�u{���uz���FI ���~5R~�� �~
������s��׎،"B!Ѡ1&X�;�iX�ڪ��[�;_��tEyz��N��L(|�~������*6���W/8a�J�Q)�I��r�ߵ'ƛ�i�;������eY��n����gv_��ZD�dK�Lni�I�$e#�����!\ˌ��b��\��?�ift	_w�^�!]�b��&�5�1
�j�#{�>-��a���+WiϷ��R��K�9��	��gwY 0H;�[{��)�7p��*}�Q`ڈƅ�3�M�ÿ��9(>�2
��Qp'�]���X+�=����̈́}����!�́�@9���?RY#x�\Cf˞*UEy�6(��&���ŔH�LkH�17h����&�3'��:Jz�Pq�`�V.'������o7��Bâ�W���n^Wy\k��'g���T��k�˕`(k9����W�����=f�=M�wO�)�Ȭ��7�&��G�m�#���E=�V+MĎ�������AXr@�w�'�q8e��C�U�D����@�0��X�_f������`4�͵p���b��+YP���O`^{.x3-�膨��@�tpo����^���,�*�6ɻ��Yʤv��E����b(�fX'�W̕η�O�O��]����r�q[*���jW����C4	�ݓZ[~x׵�f��f��gh~s�e��w֓��O��T(���;cdF]��a���A���'�l;����^,3�|D�3��x��aU�:��Pa.R
�B�=��� ��2�.b����L�R��uS��W�vW�i��nl��0;k�٪�sBM�+�6�^�d$�
�k���}�w"��좳�@�ne	�۫۟*�r5_�rt������
����u�� ��N��P�	���+c�u�a�G+ Oy�Ι��[@N����ݒM�R��@�y� ����Pr��)N�-3/��8���?#;?_7��3mK/.P���f��ԧ�3e�iXn����V�`h`]5Ӗ7����mM�/e�f�9�R�)��o��%�2��qH����a�E�ەI�*��!of�.Q�{�X�e�G�辯Y�C����N�J��H������BI���%rT� ;*�Z� �������Ǐ�XE�R�(xP%�s}[��RCp�WL!b?��;��E?�J%�O�t3�����i�����j-��	���E���fK�>l��ў���h{;yGdp�=DY*x�:�O��P$\�2����8Pd���mKv�CBa~T��5��U��\�dm(� �>���<�?�~�$>���<'� �UZ����=���\�݃<�˕k����+=q]⃡�Jh�2�[��LV_�𧻓���	�p��l?[��i�}�H�+�����0t>���4?���(g��rs��[lހ�X|l�,"��M�D�W�oYj��b�w����h�_v��7��5�n�jQ�K�n�d��(P��ǩ�2������VW��@8�
]Rk{%$ԙt��ѿ��y��2���%�o�'��x���2�XN�%|3���N!�^^��7Ҕ{���;dU��!�����?�:I���(>o��I�T.sd����|�}X�g��vd����� �C�C��t1�zը�)��m�ye��MU#��$6���E4�p�L��^�����(<�_���,�L�A/�(QlX-�0zy�?|��"̲���j�L�,(d���LJL�}�uY��v�؟����}��ɾ!���e�rk�A`x��x�ؒ�&vI��s�<�����c��s)�ڶ�<<n�s���iN�\�<�W���F���|�&@�<�F5�7����*��R�k�BX��{mMt���@B����|`<��?�x(.��뢬�Я\[4����rP��7�}CX����b"�$w�^�X��󱉶)��i�u�6��&��6`rPؼD�/��;þ���M0�E��D���Ն��it��e���cJ#�2C�����鞘N5�4��\Ⱥ��v̜��N���s��,2CQ�Y>N5��B=���[�p��ŏ�������2ŏ}D)7�)r��J��ӽm�4	fW��j�A5�q�=�" ��F<X/2rB����e�����/�]��$M.X��M�J@SW�En�{gP�~I�7�!D�ϟ�~�S�&��.��c��+�4��E|U\��)]7b	B5z���S�:9���U���9���[������7`q�ho��v�>�@�!����9r;R����)l4����o�QҒfn|ơ�/}6����I�~��]���*WN[$����ݢ3�StմG�:9�Q577T��$�)tjX@��A�ڭ�f"�CVŁR��^<�l>�"k¹8;��Q�f@��3ep�rzTm�����1��x�8�YH}4��+a�,�+�	��n,��?�7e==W��f?"�������[`��AF�@6��n��A��C/>�4�9 v��P:0'�����=J��%"�E/a����Y1$��{�@#���7(P1�䞙�\!X���SG�܆G�p|���lD���Cj��Yz����!W�~�/"9��W7�0@01�j�����8'0�`�Χ�,!�P!2O��$,����o�'��1 ��6�¬6i��ăbZ������T u�<x���y��-��&r�R�Pu�C�W�ˮ��$I2-鍩y�6N��B���b�A]-�׮���֍��ET�6�t�b��7Լ���k���	����j��7/���;a�E�B�6W���ZO*V��b���2�~��u8�ŕ�v�T��e��a�Rgn��5%�[��v��HU�E��OW�Qg��7��C�c���k����4e��:8%^2~