��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���QΠ�F�p��������m܇�+�˺7�)H!A)=8N���`'��N���K"��}�m�X��J� �e}�<���]���*`�F�Y�EF�9�j�ChT�1_ ��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �& ����*�Pk���<�T2���݉�a��<�B�t�7$@�}��K#L!9p��ud��^ڵ�@j��Ff{�緄��@~�z���G*FIC�����J�S0��
j�xp�M�,���*�rBQ�f�7�d>`��i�˄V��#0� )܇D��*,�J��p���@奈6����o��!K���ռj_��`+Xf�sO�o7in��ۤ��C��6�)^�ն)�Q����%���&5bn��~��M�c�=t�ָ����vh �1�Ъ8mS#XڄC��OV
�eKXZ�
��A��c$S����.���p`�w>�	�_	�< P�y1��䁡�<�?�(\i�N�R@Y(� �~��;&��*j�"��l����t�E|��w������y�;�d/*�D����C�34�I����`L��7�Z����1PZP#"O��ޗi'k��a�LX��9�_>��Y��o"��s��xT��� �I�P��7.���?���2� �Aι��Gr^yi`�h2�P��-<bZ�����梌��,�r��.�|��,��g�(܌�$�r߉;�e 
t�6� ��V91���:`]5v�$}c�ƀ���w��.�_ ����Eg�u�sl��&o�e��1S:?���uD�@Νt�.\�7��<�.�Y�ڝ�m$�a�,ş�Җw�!�_�n!Z���h|-M<�9�� r>�,� r��o�{�(E6���� ~)���<%F3ٓ�����
2�c��e�vםϸ�>ΈA��]���?}z)��΍Ρ�5���.�fIڑ�Bܫ�]^��Ta/pךyy�V(�@t#���,t�B�w�G�塁����4�=8��ft�a�V�Y�sV.O@3xLKj��Ê���A��xW������{� ��yf����'�ܶ-&4���57X�,��Gp�Ф�c�a��4]�9c,�d��ВG�H����[�Yj��z��ϐ�#(F�Ø�����Y��DA��?G�0
W��W}\�
+�_|������3f�0�Lhʛ�dʲ�#ݵk8������;���k�Ƶ*2CA���*I�j�:���������m�.��|�t��35���}�����>n�:-=dDH�̘�\y[s��Z��n5�?����<e ��� [jx*XN�%��
����m�RŉG�^B�q$���j���L'M)���4.������2��H�1�D�lE�����i��
��4���hЅ�+�����>��9��HLv�t}Qm���H���B��-]�f3��-� ,Y��Xؤ�|��Tc��k��������{鈸q �ǝ��~���E�w�G}\bUWw�b�펐	������o$WT1�~���I�d�%"�9��t��3�y���H���;�"�م��f�� ��b�5�y�^���a:/�n���lΝD���rmF�� �n�S�~c)��&�.:M��BFPI�ĸ��������UE�`�������Q�.�;��O*A$T�P�ޔ�ai���,�A%!��â��V�lm H��*�a��OP�˪��Ӑ�@��TC�����+4)�.bL,!妧�o�4'��	9Lk$��XA}�>��|c����"as4���DѨ4a@C������Q�=I� 2 �b.��ƿb3Z���'悺�0;h�h'����cYҥ�k5	�T"@�P���ԏ�_� m�ޟN�����D��X��#3.�T�	b�8���_�)āaD��B�
����a��
Y�hRkF�"�gL;�}�ϛ���PP+S����� ����i��R�Wq?7d�3�3���$�'U�⼘���� �?V�ZJz�G-m����c.�f�\���Ps_�o� �Jo:mi�,�j;�˜�H�%<��H#�.���mZ�k��B�g6,$'��I��ϧc���`��#Ҹ7q(��q��>��`��su5���x߆<�d9-���;�mՏ3O��y=rM�����R���D��'#��y�eM�W�2�~D����z���\<���.�ҩ�#O.�⏓�{�mYqߠ��#��@�r�&	���A���)���H+�����A��
T���U�`�y���$ ���ot��#��\ TGs9�=}�"d8�L��?MzE�:Ea���ߧ�*��_4�Fi?Ԗ��Q��;�.
*� r���la����.��bb�J�5Gڱ��H���qEN���m{��&�t&x�Z���{�	�e�����0�E�����w�<ґ{�;vd�����7�Sх�(�7�:���ۍm��J��<�e^���D2Tk������H��)����}tn��'8���6I��{P9��=�'���|�]�a3~�5�$<�4<Z�R��#ܹ"� ��ѿ� ����L���~2���1���L-&����k�v�I���u� ���&Z���+�4'���"m�G?��(�w�X����L����0�vPky����;`��fy�X��:�����9b+���*���8�8� W�q:�Α�~�"���C�cux9xd	s�Y\�tS�(|�솕�A�B��x�v�z�M�cC��݊g2�FD��юG�?u��,=aU"3.e,4�߫����Ð��i9N���p}���b|���{7`��Q5� ���o�����Ӑ��e\qq�Y"�]*�=c��B��S�N����RT�`h��!���<<�PNLr3l���h�|Tq���8��a��Y����}�Lx bS��X��'�T�x��u���kaf a�V=�.,閇��^���)�.ز>t/���R)4�L��d�M��@m�F!G`�t�����Z�%���ç���W�¶M�O�fjg��Cm��J��ѻx5L�8�yz���)��� �����3>l�W��X>��a��m=�CtZ���6�@P��
���j6~��w����$�ŭ�̷t,s��ʀ��N3����@G�g. ��׃ c����h�\�[�g���@���>��P�;!9��F�0~�p�z��9@�<��BO���9�&9��"��fE``4A��v�W�p]��K*�� ����%J�EZ9��*����/�n����ף̒��֢��^'�[�5x��}Z�+1�%-)��ѸGt��/�z��U�Q-K;Bk�7����\���/�{Ƶr���P@����1���>��BW�[��"(Z�ދCc���A��xzK�`�Ş�#��MA�������pT�x�P�w!�'Pw2
���DDq�7�w�\�\(]r�}�H��� �������)J�/�� �B�L̲N�1�e�1�S�cߺ3H�#�d��KQФ�d1s�ؠ��� >�p)�C�j�b�X���K�+On�yZ�V�< ���)�vqI}�ӱ��+Hwp"d0�yo�F��9�Iӌ@P�2O�y� Y����w�I:�����'���j�R�X�Ň�c��z��s'�Nx���;C��lG�gX��.�� 2\�+��#������y[�y�b��8�|}i�`sTP���!Ȯ��m��M�:�iO�@\qb�}A��nRbM��k:&,�	Ӱh��������@l�.掜d��9Bz������Fn�W��}�z��sf����@#g����|s�~N�������wVM�&;^�Oz(������Ew�Vd!<����sj��O�P�p`xV��&b{@R*k��K�v�.2���kOO�ܵ���$]��ϖ��EQKր��0���`-��U}y����Vp�@�eF&�J��l��VڋTH"��G�р�<qYP2F��1M�Q�E9���y��WC����m�:%0@љ#�O��Q����d�6�r���*�4����HS�n�~�sY���,��pĒ��_�ֈB��T}�������ૅ����=�Vub���WR\����_�Nx��nwM����9�KQ*u�"��@ .�����x`���@#D_H��h���"�Sr>0�_DYn�}�j[]�ڒ�a&h�F@bF1?�w���6��A�)V��F���`�!?����"�Cq��!��@�m�7�������PzZ��@B?<D��'��nɌR�b��H��'�ThYD����x��Q���b��0�E�XPD��D����%5Y'د�D/ �F3 ��D�����c�X�sѧժ�r��߭�GF/�B�?��1+a,$�.��i��}�)x�R��_/�;q%���/+�0A��aa��^ ����`Dn2����-o��i�;��g~�Ɠ���V7-2A�7�'��9(�0���0%~H�<���+��ݎ4ZQ%���Q(b���o~�_0�j�8�K��b��8*T+��ڢg�F8����zu�/�M��o4�8��s FݙB���R��<���e��5�G9H17q�%��@z�b��)	o>y����Y��35��9�i��m���G
���Lο�z~�G~k�$>p����H���	�ˤ�\!F�����BUH�1��4�X+VFw.l|�A�Tc��iQ
:�y�3]�����Z����~U�L��WV�3|�)��[暙[��o��G�CV;�B`�)���&8	L�Ka 	#쫳w�T�F��6�<�T%��ߚ���:^�	�ӳa�#Z0c����I���$K�*�V5��H��8���`R1m�^��r�#����%U�D|�N[�ꈊ�O�`G�p��H~Ҟ41��{3�)�9��L(p�ǡ���tM�'5YC�Yf	T�'��Et�9lR{����`��)���Ev�j�[�Gî`x��K����x�
�E��s��K�8�-���b�{����tTI�ܟ��#��=o�AEߧ8ccs��������"�n�:g[�.���f��~^&��p)I�����j�S	�w�ZN��'9�@�����JrQ�]i
lfy1%� ���)cㅲ6G�G��yG>hA�g�@��`�3�@.��*u�@���8.ۀ?aL�or���>��vq&?a���_
�r��Re(�Cj���E����F�z���ƈ�'��Lp(\�Z�&��P��d�h�!��'@�i��-_u���{VwL�%����Z}82o�PA��6��%:�c���J}Q�OaT�uOW}-�W�xSJ�I���H�i��43ٯ�����u�,��}�Sf��p�X�H��&��O�m�Gs���]��ϫ����Z>*��������|>¦�����F�jZm���)���qI�Ex�=5&���K{�S�b �Z�X�2\co�A��U�G���*�8�d�w!ч�À(ϳ�W>^�U��I�F�]J��`	 Җm�]�H6��1��%����s�T��6��~~>;�2V��4O4�ov[��"X�8��.�E�#P��7*�w��M�v�`�Hu�畊5	P���a���~h=X��Y������������Z$�9GV���Ȗ�X�ɗ�v�\Lu�J���"���vʷ����0yuQߟ/�� H���U�n�W4cଽ�� 
�Y��ǅvә9��w��`�O��g�v�^��[��ٙ@v�w��^�ey���uJI�A`�,%� ��g���9��WݳM\�����`iq��'�K�>p�Cm'y��zS����u�w�,�����s�'�`�ݍ��ُ /Dƒ�P"���b%_??�D�e��$?�&��w�-*���M޵8�W�����������<qE�g|1�7ܱ�f ��jH�'��oWG,n��R�Y4/g�3�Y_ܥ��)$m	s��Zm0�79d�M�]�C�s�3�%$(]-�'�9��+q2�!t*�}�H����֢��S!,E�$T�E��@����]O������!��^�v�t�̃�Z�@��סq}5NT�~z{��Kj�"�"�	�\7<wu�7m�Ni�h�g�ҟ�+M��0��a��c�����ʥC��?��C�悆k�J�����M?�&�g&��$;+�t���)�2�Ɲ��r�؍�T)��@��]�a�A�	f#�@"����܄{G�w��4U������Ʀ7�	|xCcNg/_I"n��e:Gy=|l�����T,�RZ��q�m�5ْWc���&���� ֲE�΢��ڊ���']&��x
�n����l�Ң�%�#��چ���K��]���̠$^�Vz��4��N��\I��;jMGk������5V����������]�ٱf�����M��A]+r}�u�{���$f�Gq��)���*�W��lJ%4Wv(��*]Sh@6���gY<{��o�m��� �#��`�g�$\Tw��u��n���!�s����L������r� �Z+�����h��赤#A.�CCH˕�?��G�ٓs�/�Q���̧b/����2m�#�6�bLDF��L���T���_�s��:��U!� ���3S�-���'G�3*2Z����-!���E-l���Xd��V�����㹫��26�G˓�����0ۡVl�Px��7���f�?$�D�l"�i���.�0W�h�i�Iے����,�c��T�8ј���������,�ah� 8�L���"^���]�0�.U �.�*��_$�v� E��d*�CjH(o���E��͠.Dm�i,��m��P�Y@|�&�uM��}�\��и��QhӲ�b�R<�>��Є~]
�j���,gv���&�����E6�K��O��lZ5�2�|&��Y,7q7��D��u�K��o�v�՞�M#���%���J�ZP���
O��)�i�6_�9�C:��W[l-����z�F��P)�[Ia��P�\qjw�Z�Θ=ߚ��1����s)�{t�̛��Y=���*R5�M��T�`�(i��&�;����5��O-�}�4m�4���
�\�>�"D�v���k��7x��?���@Ț�:�&���U�r8��H��%�}��:͏�dY�]i����t��UDwL$~>؎�g��i��ئԒfY1�l�+0���߾Q3'��H������?Y�ҳ��B����d*�5���,Ar{\�u�t��h.��q����I����y_����f��Y��Ҏ�$�2Q!Z��qD�����e-
wX�M[s�J��y�T>�p���Sv�R�]��*o���l��2Z��e���@� �K����0�1��!�L���N���}b1ܕ7�������7'�L��V�55��i[()����	_b�%�v¥�O8�(X�>p�lc?��1�C�D��En�[�?v%c�Xr�=C9�pG�� ��R�[��X�Ŷf��j�O�L��"��h��-�Au`ܕ����޵�u5��v�XoAWE��#�ǡ�p\)v���3�B{'l�{e�ʼ�����q��D��e���$N&��X~��X͖!����Z�S�ڛaKN�}d=��
E�1�l�ٚXY�>;�bū#��Ge�3���SVI�
�O,��u/��ϵ�E�vmj�V��
�]M� �Nj�,�k�܉��7�;����P��91)��p+�Qc�"�\E�bӀ��>��.�Y�ph��L�n7Re&
?8�W��~���D�-�[���r��������"�[K�~���}��uJk&�ߋHX�����|�5.�i��3�&F߀\�����΂O3v;~�7����ϨϘ$Ow�Z�=��Z�z�0���;�o}Sy�U�2� ��xt-�x�Nz/��C���o��k���2��oxi���n��%�L"��P`dsX�;#�#E��X�V$yl'�@*�Bs;��c����oFj��K����8�|K�Z�k�a1J����4A���X
w���@UBQ�[�@��]ϳ����cK��7d����q�#���h�]B�~�ח�s��P�r�`Q�]X)�$jO�����1�e�8��Ã w[�M,�ޠu�I�3����^y=)�� ߆�H�4��}��������S��Q�ba.i�I1�����X8+h���H�c�%r�wK���߁�3L�*ל���*)��N�vO�����W�MP5�i��&QIX	e����_}�Bq��h4	��m����Y��뤪̡5��E{&�.��⾫���O��2���84���S�(8t5阝��`��\���s�|��L npm�p[QʄàWdI[��t1�p�A[�hs��.�9g����*�sΕ�j�.���-�2!���$0_jd$|u��I��Q�b��'k�o#=�b4WV�S�| �019Q6ۜ���^�4/�;�Z�ł¸��z�m��ۮы^�� `�`�Uo��?�xH'����ۤ�v��ʰ�(��1OC[K3�r༝��(���fI��G��4������n����G���3:�NĬ�민̏%z��J��G��̗�$focM{%@��_����k�<��x�H�I{�Q ����l��AE@�y�Xbb3\U�H�?΅���ڰ�����2��2o�
lI:5���T�b��{�N�=��<_�o�P�X��Bt_sJ8�3����i����|F�Աi̭��j�eą�����3���'_�6�S�sM���$�f�>��$&��WV�J	wSm	 �Y;�VV�r�[j#�m98z�F�����L�isN��Z3w��$A`<k�|d��uW@��F����I���L�a��}�#�R��Rf�_T������%�K�\��FX�v��[҄- ��An��Z�±�ӟcT���[�T"�k�X�v��T����ņ
�|G���hϫ��|�eʝ���~���|�:f3?�U�))��.<�*��MWG%\�aK��m����GZ��%�����8��M_�ю��cO]��h^��A��j?F�a	�¥���V�bϖpa��xp֗��d������_�V��jƃE��%$��A��H����N[�PK�w� ��a���\R$'ܣ�z�)v9��8W�Z���E]M]P2/�!{����q�Y�
��R�&W�9h�"���Aw�*q�|�!�"����v5���:Qu�f�#�l�p���E��֗� F �;�:x�Q��.L��?�$f��c9T��
�����jh����P�hw`����`ϼrwe������W��e����a
i�zQN8�
S��)-*����`�+`�-��u�v����r�=�񊓝�'` =t�-�?I�����Q\U�=���_��A�1
n����7b�&�u*�y��S!H�f3ϑT���=s��W��;�`�&�E��I�t�W���/w��5[���a����"j�r���\���"�����k ���#k�-��pU�'�'�!ܯ�'%Tt�c�V���t��oҲ���٪������w���&>MK�5mk$o��S 0�X���cǴE���Y0Y��v�QHW� 8�q0�|��g�\rTFܐ� ����JB�8��G���י��/�O��,��]q�D��)C�D����6g�v��	�:f���c�[Iem;Z׎�~�R6:�t(X�a�kW�98����e~VM�FO"v��mIG��0��Y=�;���s:X]�b��:�)K	��ď�^�#�V�1V�������Xܤ~����U��x������O��%��VFˡ�Ș��.4b;��ƽ7�3�ֈ�E�t��-k3T%��?��Ϧ�LE��+�������-�a/��9ߙ���$`��:O�+'	�(g�F��M��͝��2,������UI�NݒwG�pl�*���&ڛ��a���#��v�ۙ�~wW�b$��Y����z:�~��������ج����_L!Ā n(�w�.?�N�5��bN	
�m��a}hH�����ԋ-R����Q�^5Lو�	3{�ذ��)�B�_�9܄�1Z
�C����]���u�1[�v�۝k��&	�5y'�aj�n_��#�G��ۘ��X�|ǀ1S�OY�aU-�w�/�(=Y�|��Ga^��D�X� ̑��(X�׃�i�Y~�o���f: T]��ģ��8�F"w��@ܰ�ݙ��:�����L"*Tdp07Yҋ��]�iˡ	F���T-Y�����Ȭ�h(ԦSMh�fc0�l�r��_}�ξ��ٴ�.YD���j�b�(Z8=��;�-������S�̌Aė$4���bz��1�ȍ�Ŝ���W����������-`b�p�h:o!�����q���J��Q��F��v-��7>�� �̭�-�Cl�l���bn[XB�`��Wy{��2%�@�UM���(�o���a%�ꭍ��K��;d�o~#Zvw�g� Iw�i�h7#��"A�Cb�;��!���ۦ�X�-uE��K����9k4����<��τ�0��+	�Be����D'��ţ!����`�Eti�j�兖U+���g��m����މ�_K�P��" ��"� ��� �?�w�aj�������>���g��:�$���*S����~iqx߇	�L>�|�t��fȠSŲ[;vwW��aSS�mz�E6�Ǖ'.���"�p�;�1W�i�[W�_όe�ihu��j28ռ?�Q�?r�`��9�B�yI�����\3�z��_���7S�y�7�Hk�r���H��T��~�|N[��1��4���N�#�&��ܭ�ɐ����#$Մ��Q
5��ӿy��^�˸x�>�PA"�T�
��&��Ⱦ�S(Y�S�,�����)w&<]�u���3��Jt4=w���V.���^��W6�G�N�ۍu���sN�!�N|h��-ʘ��tRJ���Tv�i�M�&A�xK]}�)��$�A�V�M\uxS����$�Sw���`���m+(�u�l�B�WK�\"��� ���+�"_/x{�ߜ�{:����J �/5���V��������H�C�g��kI����
+X5�=	�o�ڰt�I��G���_ ���4��Mg�)\{��Ҋ��4�����CF�k����t]�ȕ��yŗ�@[�L�8�HT�96�M�$���j����s�Km���@G`��I�ڇoήf�k�s�Q�0�Uky�⏮5h����M��RU/�g�u#�y@Z�|��GX�����9���z���>� ��o�r���l���a��)��d1�&�o���\���i�������V'�GB=�Ÿ�m�Ll��:�ߋ��J�)�m�\�f��e�.��<� ���7�Kn`�)/m˱� w�Nh^�sK�G����Y��.���6��&N�!��2'ӳ��U�g�?&m��w�A���v:W&�	����kՍ�@����7��ݝϧ�Q��;�B
�c26G�[ܾ��9���߽��<�G6/��!��L�����T�:�����vV�`�ζ���+�5@�{���F�E�o)L�%9K�(jĽ�AȽ�T��=r���Ws����|��79�gU�5+�=�r���R4��R�!��DZ��W+d�a���0�Yڄ2�2��&��+��ӑZ�@0�!0"}
�4��ˢp[fK�+-�0}v�����ۃTKg��Y#���6ٻ�y'�qzT-Q�C�9^�6��� �ϵ����_q���N�2�/��U� 7��;l���#:R�u�x����K�?*�<��!P�d-��6{���;�� ��z���$��/�K��e�?��<n��%��҂_R��y%d;=�����;��l;��
F]�i��-���3W9h�kk��������!E�.��`}�Z=W�$�!��߲������zA͚���@/�@�3�vi������%�R��O�P����V���161$$<���$K�L�*=W���=�9��`�T(w\�QQ���73�d�'�G��,��2fb|�ͱp�)��d�o�a�R��c�����	y�t� ܗ:��xyT&�8Me�NePĢ� {6~�Q�/�Z�G���퀚qM=6�1t��q�͵�'���У��3s�e��	�z�r��ٷ��1�.ID���}|7��ÕrVm-��Y6(@�q�WQ)f0�����>��4B��7T��A��v"�T���L�
CfD ��Ԍ��>z\����}	�Q��M�4����Xr�w�k��K����{SQ��
9P��k�L�4�6!i��ܙ���,����ۻ]�኷��T� ��xX��A1!D��
$X���x��:�B��j��"��*�F�ê7�`s}_����P��D�����x+��4~�ki�����؎��T+��Z&�L(��j�,�o=�i����$�{t�}�I�$Ԟz��?b����{�&�3h%r{f9C$���R���~/�6i��%�h�a^K�ԕ��׀�Bxh��M�-�*F[7g��1S�z�A8Tt�5�F�G���0��u�ݿ���J��}3kv��kJe%:?��Z�3<!b���r��O����M���%�rC����%�3IC�Ԋ��L�!�s:=���`��᷵�^:|��Mp��\�EK�qHS���u�F�mf9�|�R�U��6��iD�乣� �\jr����~�j�@��@i�(���y K�.���R�Q>�iUO"~���	[iI+�*�y+9�J���c�-%G������$�Q�E?�H�Eie�H�P�9w��@+�T"�">)��2�<_d<�c(UL�$=6l.2���x��l�bͺ��=����'s�"��eG@�R�:�{ӄ�!�W�E6�1�%��������ǵ���,ҷn��Im3C,k�C�`hM)�
D���z,VA�j�&1fݟ~�(K������'��μ��+��&Y��%4ߤ��=aj@II�� �T���3��jhKO�1ZL�$�>�ɮ�����_؂=&��Έ<��է�ңLS,���pOxI������M��i�zo��?\.���uHBӽ)�=9�q����
ui4�] �&j�����m+v���*0`7�����#�,Ո�b�@f�s!�VE��Z� ]����\��1�3�A��¯��pI��~����r�ԣ�0��*�ݳ�r?�7;�*���jq�H��7�6��֛�=뛐G�	DD�u-�wt`_�<=�xJ����Y�e��� Ra������s Ef˾@=f�����`61����I-ʔ���k�T�c�dY8�V�w��BQ|�pM�i��x�
`8��X�x�U��Ρ*y[4Eu<6+un���\����R���*���?I�6�j�0Q0Rِ?o�=��b҅A�.�`�ǚ�.��h��c��H��^>Ax3ݚ�I .@J9�gHF{��f�1��=D��h��kv���{��-i<�I��C��3�V�"=�����x�7�� ƚ�v�6�A���՛ �7��<��v�k�<���? ���83l��`��[�-��OtV������jÔ\:�zĚ��E��f�-��i�g��T��,��s-s�)O���|�Ǯ�d4�!�8ǹ�^����O���v��nq��:��fO�ߩ%�a��{���Ȼ���N��v�n�܇%4�!p�
�]vJ��cWihNgq"��˜`(>���Lh�ps�r$(�jJ�y8�4����,���^�)�j�BC*�֎�ـ,+��v:��n���t?Pi�W|a �t�v��$/g���|��+N4�k�nz���M¬H�|��\H�i%H��29�a+��&����j�$%@��������:
}�)[`����X5����@�{�To�w�m�mOO6x�s*��Uh�v�A�LW�CG7�KӶk9�8"!��i����ʁ(�Q�݌$.Q�@e��K䂻AD�;�7d����.���_�Xi/Ֆ&b�r	�mÛʤ�c^&����BN1%H��>��/J^>ŧ�aڕ�
`~��Fm�#_��((��溝'�pD�p7(/�����dkۤ��AS��V�箉=���z��%O���b�Taok�"TL��l�z��yG�
[<������.z��̑b���v�"���	ZL��p���������,�zk�xYI���NeWp��g:�#~K�3ʇ
�	�O��N��{\qtoؼE�)���d�GN�~����7�M����t��N����d�n��˓&Q��6� 1%Ha��e|� ��	;9oѦ�1K/XŰ�6��}�p*�^G�L*�zJ��>W��x��7j]�
�4xP�b㛈�C��X��SE`u��2l���)���kߌ�X4�ϣ$�	��p�:ؚ��p���Gԁ�J��X��Sｨ�7y�ŽųqF��z��W�)�.�qMhΌS�7;�,>c�m�Ԇ��R�~�&�����څ�	_B���RF}b���ޫ�Pl,���K��	���Jw�Q48���JɊz�������������a����!"�2�`��`X�(V�:S���7}�'Ci�?Pg�jx�6�Gn���¹m����A�㭀�����L�5a�F�:��!Q�w&����ˮ=?�%�Gn�u�Dd5P�M�Ε�!�ouX������'�$���k�*j � 9!)L��Tǋ@��1��=~��d-����v+��I���Γ��dH���:��F6p���m���cT=cE��7x{U�>,���(�Cͱ�"���,$�N _�����X/�t�)O����T�ie�&��ZM��5LRB�(�Ve�b{�.������~��y�'�l��!��I��r##��P5a{�6P�����qf�"�����-'�w&h\�n�V?p~��Q�����G?9�����7����J�X0����	W�Ҷ�'����9��D�{2[��(U6 ��kue32'�יL�]�\��t���5�۸�k�CxY�
�H�CpU��Cf�j�[C�]�{�PՂ�b���p��,�wm�[����(�ښ���V�fa��n�/��@!Jj�w�5��'([��5Msxy9���Û��z����1fT��d� ����
x[0��#7�Q�t��-�1>�1���Z\zy��
�c�G{��tE��=��p�����q�d>E�1㷛Z�����p�$���SW�zB0��� �;�=;g$O�g�����CE��Go߄Ek�-dD*����i�}�Ȋ&dC��W��Tn$u�y����3>����Tp[q4��������j�O�#�?b ��"�������"辏�<
'J[G"&�ӛ8��T>�>wE��]_�1 ��x�ݞ�v9%�k$�0�j��� ��Gp�;�E/^���S�|��r����h�վŠa�R1�
Ro�����|�8���6|�ov��NP�F�+��b[`�#D�apH^��%��m�[�����I�B忯[�T����mx4@,H"<��[�j*H�� ������(W�a��	�]�3�Spf��ӆ]Y������u����I���Y��B���fy��4i1��s'u��V)(�F��Y�$��7T9%|�y��x''p�_ ��m
((��I�,3��>U'_�����6Ǐ;=4�q�Sg\tGG��V�������,�i�\�W�O�O*]�o�ŷc�G�q����Kc�	;	�;�H]#{d4/�]���O�h�D�[��a92M���d�;��f��N�A�<����Y8G��X")ֻw�����K(*�ʧ�"(��?�Ұ��D?�^�>K�wn�jO�W*����کȳ���5P�����z����º�����|�ϣ�78L�s�jrX�mŭ[9�����\�6�d$~|ѣ�y)Y#Nj�-���x�'�8�zC���T5��W�b2���@������A4	�*�34�9N��㙼���B���A%gu�g�x|O,���tt�d��։�H��2%�>/�FY�H����ߎ�ۨ�/HC��%N<"����WQL~��)��=C^>E.�*�q���b=(;�U�c��(،��X(��00�)o���Ŕ72����	|mׁ�"�6Y)7$��5P�l�ٷ7�}e%�V-�џ�b3����"�м#�|O|X��D,��"�3&+�zik�
&�6���Zz�gz/�Y�*���:"�z���7�L������ ��!K3f!������T�/ʸ1�$�I,�vq% ��I�,�z��q�C'����9's�����E��n��7�- ��4H��犲�nY���C��^߈0�3�h�Y4�L��x�M��'5�`r�1+R^rBsu?�&<�}��^x��W�=P`St�=V���eܤ�ϧ&|vM��$��I���,����1�Nra��7R1Xt[cnC~�nTrO�ga�����ޤ V�� ��^!�iҡ���y��R�=� 	�����܏N�9W���i��E�����"��g��f��G���󅧪��N�g�2��#{��/ïc�������ވHHчe���S�M�o"�D2\A�����bs�TEp�)q:'A}����ⴉ�^�;�~l^��MC�{�|�u���w���@1ؿ}�0D��,lL��������:��s��+����cc�)��&&m}0��2~ZI���7
]{���U2���6<YW
M/`	�l��O����)�DD�	\�����,#��g �VMn����U�d:}D��:X�Er�l4�p�Td�'r�������f3 S�5��ja=>AQ���i`��N����ZPA�Z��֗�+����� RX������g��A�ٜ?�����@*���?৵�l�$-����8Ӿ�j���~�ܨ�垗���È���un���`PH)y��6U�!��b9I��B���A�}�u�9X�� �"�{a�V�L��\^TIo@�6Y#�a�^�>e�#M�G �k�jI�޲�H%j)\��xc�}H?,!��㞹\W#�;w=�Lz���_	��n�L�9#D��M��oB,�L\�u1�?j;�<S�U��Tإ�n�:`�_�O�����'��$<��%/΃����D,d�Ɇ=���4 ��#?�p��ٸ,��JV��q9[��ez��:eʮZ!�`��/�*��O|��&��=�6�y�w��M��}�8����Nf4.l�P�m���#�7�Ķ���w��gD��*lr�z�/�Y�=�c��{�	�OO����Ucb���q)����SF���9���aB:0�`����OF@�!�r(L�U؃����k����I� ���k�'�uo�%���\���ﮇ��h� =�����V��eA~K��a�,ʷO)֧�#�X	ݰ�h5���iJ ���5���[
.���AN]���.��*F;Pw6�����	|�r���#��������DLaw���
�R�h50�)��P�Gˏ�����G/Z5�@��|c��mG�����Tp��ۿ�t�P!4�$�F[��A*�0x�����@ا��湂��U`�>��L�b��B#��C�+d�d��M�p���	M�I�]�#�ǰ~�?B*�{͔<Pk{!�q΋��0�0-ɩ�J����KK%�n�q�V���x5\:ɫzk���21A��}s9�NF셳��+a�U!�7�� ��U���ڀݐJ����3Ք��4�ޭ|UH5G��֎B.���ڋE{��0�=!K�
c(1��(,deih韅]g�v�o�1P�g�!#.�dŘY�	��^ަf-kJ�=$�MVK옇]+JϽ{m���AA��V��F�&΋/Y��\����o�D����,�������Ju��X�e��;�hm��f+%��z�s3w4 2
��������}5C4�����b�7���8dM�.�D:�IࢯH�l��jeN?��ʻ�ޙH���n�޶�i�IcS
p�6��`G�GtG�W�-h&�����I�^>�p,T�=�9���0-I��p_��i	d�內c�KK$�$g1��N�Ed�Sr�n��|B!e��M6�4��ә:W����&�3s����8P�>�+]\�b)���6�j�Ӧ&cl�A_�L�,�m{<��D��`�UR
���?T%�s�ȺK��<�]�j?C
����4d)ᒧ��/�����C�q�,�z�?�6,�5�*��Ox���J���E\���V��[R�H��	��F:�(p��|l6#<�#љ}�ʴ9�0vss��	}��$0Ǖf����2���o����b��G�U��3����m�F`p�����Y�WO�۲�)s�~��a�[�W�ϼgq�n>��&R N��K�Ub��j����F[9�~�����n��]!���F>Y���a��0W��	PNn�`���	�3��凕R��_+�����p���'��aI$.�ixو˞F�Ó/63��!]4�`0�)I�>*�C�>��)��&� �
�L?Vu͖�"����2ΌsD�>@��;��0ؔ���f_ֽ�%?����v!���9�Wz��a�-�y�I�?Lb#[7k�pI�	k T�3ŧY���?ە�&g�֨��UcV�)��t���Ba��L,�~�U2I�������<U���[���q�"�iCa�m�%=�`����g#Z �Eh�2n�NtM_e���v�x�����u�O}AF\8Ig���R�Lɤqt4���u"������p���AZ�}�t	JZ�r2:�� ㌪LR��/��=�ī{f�{�c|YszUƽ_�[�mG���0{zV�$���S����e\315���Y��"�rK� S�&����5�Y�h7�-���hg��ݧ;�|B6Y�z�F�e!�D��q�
4;��dD�bC�,�}�F���Ɗ�(@i!}yq��r����+�I���hh5�\ �)�r��ͧM$<�ʉ�l�i�G�?��H�W)�u�"�q���t�����e�g��+q� Ur�M�b�ŘT�9���Î+A�J�=i��/nN9�9��ȕ*��$nCPΫ.<�rV��m��/U��j��i�.��^o���G����*xs��Kg4��^�".c^3DW)�0z�1���mUz���q|cx��v�n�"l�H7����ͼG��ܿ��qx}I,s4�x��EMÏ;U��63='��8�ħ�p��h3wvB�b�4�������<��8U�HV�A9"�/Ъ�cjG�)ļl{�7|o��$rTc�g�0L7��ַ��܀�����+f藑Bm��^��'m5>��jF��������a�
���ǩUq�V
�k�M�9�:���k�^���S��"$�`R�%�ɓ���f�qX��+��ZF���19�P�ʩ��t��89
��B��Y��8��6��JO���|Noh�q���J*����[��(������
e׼�D�4'|&���A>r<)�������r�_�K벤p��Y%�L�q�����h��ߘ�Q���������
�A�E/��и8̍���ֆ�ND0��g�3�f���6\fJ;��rs��K�*�]8f5,+�Ք�c
�!��eDn^A�?X3d�t�k�+�V>ءsW���O���^A���LdɊ͓����_-���	d֒vwq�pmI�C�<&Y�/`$�kU�욓��\���ŝ�̰�����V�@2�����:�
n��>  $�� �Pz��)7����r����lO\�k�	+��u�V�`�=���R�{��:�M�5>ڨ��8'���G ~#G��eD)nRG9EA,�Զ� '����vZ�{%�����LP,H����{a��o�5�����$UGΔ��E�B����W2xG��N-�#ڠ�ˋ,2����k��%����+���z��XG"4�mS��$0�ʑ
}�E�d�0��Ь�kv �UQ���/�Su�@#�>� Y�4��]NY�ߙq0���;���fG���T]e��d��,��pg�@\Z��H��W�,���.ܨ69�{��W�����:�u�te�Y�0f�%5�O2�d�z U��vDMKmP�y�ˆ˖ͳ%�v�-;�oMY�vZl�K׼�v]ب-��7���M�>_x䠶�=��l�-:��e"��D��
v#�Am00��nҭ(t���G��������3/�Q��L�@�l3U�Z���nd,���l��2���Q�������3�2��(tі�{7g�fTP�	/){�#���	���ۑM�`���Yx2�A�n)��ds�I�W�z���kt�qL����K@�b��u��a��\��"��g���p�mNo1�a˂��\�"?VN�~��US���wo��c#��Ìs�ԝ������b��K�� ���X[҃N�XH�8E��ԡ�����͕q=^�V'ج�U�8;μ�Z����Q�!(��7��=��7V����6i��x�6��q�_C��3Y��`�5���|F1�۰�^����^����r/�wu*Ƭ#�Ń���-v���G�G3r��>�("��Ь��[6����^4b�Z��<b�鵆0/�q��T��4���j��ˉ�e�C$�2���v��pĬ#%��p���x/}9q�h��X�4 ��"��0�5q�o�5j4ĸ�Mԗ�4n4���0�w�?���emVT<��uAmI�`�R�5��Qc3"�yQ��_j�^	S[���mi�h��11.gEF/GW���Ҩ��6u�r,ƶ�^䡜���
Τt���C�eh'9��<^�Z!� ��6e��1��)�ն]��ĸ�Co���v��h!q�-é���LsT�͂Ь���(s�R�hR�ƍ�w���πO�«�Z}B$��m��b1F��ɳ�3����'h[^�?U#�w��9aۿ�4wG&r(�J��Ć�[d����ń�C ��r5�s�X��k���|�{j�H���<������0�Bb~�5�z��-Giη��!5H�n�Jn��s͙��)�d,��J�����n�-�R����zkĲ
n�"�Cdfn���c�z��d4�?�3I"��\�a���q�����QG���e��
<~j�4���_����"/�.lA$�G���7)��*s��ZITo"b.�^.��++V���N��fybO�xﳺH$ڷls����l&��������X���N!�ށ��mKj?���ZiY�;E?GZ糩Yr<��Ѳ5��O	���ݣ��fI�gBy�=��hI���4�4�%�>ؙD�q��ݦ��E��0��c��D���t��d��ڤs��/�;"���:چ7��g
���V����3D��,e��y��݊����~�7&��+�:b���S_�f�C�Q ?�2���Q�mf���t���Q�Qu�a(2�U9�aD�$໖��j���"��d�=x��u�F����i�͙"Fr��AX�Pj
n�'\��y%d.}%J�@-�)āje3�}��f���d��c�F���\�8T�<I�A�i�Uc�+��}ME�k��T<�ܩ��
�I(���l�\E^��'���v���&���xg$�����G}>���0)�^�q����@�;m᳑�������ZK��C͟�T1�x���ӷ�������WX�O�>tGj�酒8Q��*Q�,E~v����\3V���x�Ne�[���J�M�U
�t���c�r.[��U�t\�owoM��3�Mw����lq[�����B|�`�`��x\צ���ODKv������D�O}fC�t �CPDv�E$�J�0��uo��u���{*����;�A*zo��!u�(���"�y-(DP����G����u"�0D�i�^�\�+ Y�����f��&���[�gи�mc�K����K�nl��@0���>:�<�c���5�U��H���Ddԅ�E�(��@˧�l�{q�{ Y��8��m��V��P��(S�e>L���NO��4�g���cK?����}s��9{9�0+��Q�ڕM����K*��n+\��>�-��x���1�l��(��h&�+SU�D�xLg���t%����5y�+�˹�4�o�O�nct�ZQO�t~>�_\���a>Щ�u�c�8�σbC]p.�p�΂���
1���/?��kc�7E�p���K8aV�ST�+��՚z��d������fN���XN��3����2�[(YJ���_����]A	ɫP���NW����A	.,y.6�\1�z)WB�$�l�O������}������K�'�f"^t4�)*w ��_2N���F�~r���O��?ɚ�?ȯ��`����W���ߛ�c��D��m<ΐ��K���n�l���'\�^�Y��Q׉ 
G*9����+3�$lC6�j%��$�W�A����
�'v���uT����)*H��)^�a�z�`��Y�\�WP��?���F\A���*!���Y�$��<N�l�׋+���Ax�3�i��hGA�$��oë	1������=�&�5`�z)?��;�o,�"D���i?<���&a�I�Z������sh����3�:�m(nP�2��J��_�kbZ�.�
c1������5K�h����_�T�}&��o8��ʔ$Bσ.A���tKsU�b�Tx��"����guy;j[�P8�nP�T4�z�{���Y,�b����p
�i��4%��a	�FL#�)��4�
��a`�ܤ�� �%�T��+��Cih*��MY
c�0řuHUI��~q��L�P�u��e�J��n���U.6�bOf��,l�V�:|��vARRL#I���}��{�7'f�+���N�&���G��0?�\n����8�A�4l�8�T�P���w�Y��B'�0v_O7#n�Ⱥw����_4~q	G&����dh��p�c�_]=�ᰟIay�Qp.�b!oѱ�Y�gm�&煪����j��Er��G�:��y��������Z�N���,�҈���B-c��d��C������O`���ߐ�U�X^hI�d�Z@�u�>���ߐyHN�c��SU&�i�����W8	���k���U�,�G+y"� _�d��oU5)\�*I?Z�>�++gr�p ���g)^�[��ï#�2~ŨY+��"a�ߝ�A���퐒�2]ۥ�rI��������c�.A�&L���X���1ͤCT����|-rV7lc���w�g�z2�H�lUX��ݮ�2m��G�^ŋ�L���m�`�"�6Se��%v�Ď��U*ez���� wL�_�Q���z_����=�a��; ����2�47����(�?�rx;[œ�ko6���I"\9
��������Cn� �_{ߤp�b�7������7"�bd��)H��R��(�>�R���2	):xp�G�p>��q`F�"��e,T#��1MM#a�S⡇��I����Gr+m�,�v�U���a<���o�暑�5�
���|�2E`*�?k��|���R >7~�]�'G���!PɅ�g3JWT|����m�����Y� ���":���!�t�Z��e;Ô����k�` iu��EPZ���z������h�LW���J^Q�4P¨or��ם��G���� "8i��������뭵rg���_3EO��(Hg|�R]Fj��g��b�\9�.��\U>�_���%�b����g&������s�T'N�ql���DG�b��(.` ;:��5x̱{Z��X��%�˾��Ն�Ed���1��!�$]e�{Yc���{�ҩ����yR@G�X�`'8�g���N�vvo�hp�l9�V�[#��9���Û�-&d�Z={A��d|�×=uO&z�i褫�L.�"�"[�k��2����S���-i;�?Y�j�˯�̩��I�� �σ�)�w�')	��܋"�a��>�6����M�t�	n�9���?U�z����m�JP���?[��q}��d�ю`��]���"N���Ѱ�z=��Ձ8����HBw���?#KU��-�y^{�e3)�IZZ&�@��x/�\s�A- X�̚~�Xk�~�L��^r
���%7ך ~��e�G�_;[���=����l=SJEE�[��*)�]��>��8P�։�Xߨt�2�c�ж��k�
p��3�Or]K�9�-2�[P���_ t�#|+O��Q�t�u�E&�sGK�2u���Z4�%c~w���j��=�5~��jWa��q����5�غ_�rL[�p=�{,��0�W�
�߹��x���*�� :�zZn��Xμ�5{�+�Tei�v>1�ߎ:W��M�����r�W�U9�����ݗ5kuːV�r�����1��s@�4������}e�����ݩJ?��K���F�φT�OҔ�Oq�!	&q�K��C�}n'BH�&���F1j �pYіST���픽B!�/�K�jj�!�x��>�'��N�b�IX��\���P��22$�dmrT";jB�����G�X�2ѷ`BU5N��?kQ&���;�a�3vC�B�b#C-���~1��SWk�E��-p�µ�������0 #r�Ϭ|mS��3{�t�o��ǹBq� ���W�Mq|��>#z	�f!3�7�Kj�;3׊E��s{�O��w�Inym�-��Q�w���#\�F2�źB*')�jNg���#��G��G�0,i!�[Ҝ	C/Bl�(�6ϩ�+��N:*�C�m[[�!}0$����@����cb~ߝ��ȞϙPfW�l������Ey/� fKi�xwRG�7�D6�.S��q��2���R*p�{K�3��`cc6��L3[�&��i�����	��ڦ�d`��/�=#�Q_+l�������~hϾ#�צ�s���fCd�U:�q6O͗^I���;{��5��7GUv܌}�.$��%��GO�J\
�|�ɧ �'ø���%y��,����@�!Io^��QLYk!*]���-�{Io����a��xq�x���f��{[�^T�/��s�o4����������I�:䉋���1�:s���1T�/-C47�K!�O׃2qb��&ϻ��oKΟϖ3y�A �����ԫ��:�m�3���A�����e���Qb=v�������Ӣ�:C�*��:�i���ݙ�:7��S�q�GД7�>�\��g��La�ۊR�K�q�=��'�^Ú6z��BQ��0�b�a�ZP�9�";����}C����Uw<�F| �X�j[�����_(�����)e�T�rإ�i���0� :���8j���q�\���w�	��/wo���J��;����怤�8�����d=P�C�$(�k�[�(?���=MW3�.�h��4��и�b�����oA�@�����DrߏyK��U_�)Ư\���b��b�!�����P]����b���75�T~ �����=L�Z<_�;�0<����A��&z]\�J'�K,����<o�	fB�֣��$��ajvۀ(���)��4��o�c�6S�F}<DZ��7A[��*��y�E�����d�U�Z�?��M�u��Z�&s$3I(/Z	p�Ɯ �Ě(�XP�<>)�9)�ۯz���qh�Rtث��y���b��*�I�x)��@4��2��-�m^+[|�%2����G�8\�3_ ��ţr:
�4b�5aR�#��$�`��#�`ʌd�SNJFK��I�d�:��e�lo��{9�s"�{�׎[Z)a
 ���$�R���y��ZӨ_���2"W�M(8���?;��Ȑf�sՈB��r��c����n>�CVq��:�Y&��V��7p�
B�D��������T�k�(�-����+�kaܲ�6ֶIj�Cg��Mf�ó��$\;�>oD�������1��
���6ѥɥ����!Zir
���Ȏޜ�!�5������]ŝQ����B��]�������T��\ ��� ��X�`��e|̶�sOL A������\MQ�g8Gƌ,�UBGil�P��9ڌ뎺�I��/��4S�*�'w�(6�p3 r༧����J�?@	Y)Pa���2n�c	�AOrEҒ��nQOe��0"a��$�ڪ cdn��zO.-�h�}�7���̒���E����Q+u������b!���`�IdL�if����A�C���}�f? ���m4�F���Gw�q	w�v���T�$�|�ߘQ��b� T��+0��s�*���e�}�UPRۅ'��3PK�tp#7��f�]�
t�hC�������~�/}�q��xb�{ez���f}�Q%�Q�Z}~)6�i�ه�r��e&�V���PY�(3o�\<���j�,�s���3��I7�%6�ld<Q=�LgO
-"���e�������*�b����p��������I�Y�2U��hrB��@� x��ږ2KW���vS�/yd�T���먊����/�3pR �2�IȽ��>������)�G�!�ljs�N�)��@��oM	��v���͜s-$���:�'
��z����(Ќb��j�d8�X40��<�k�u��'�W0?�V��l%V�.O߿B�hIB=/W�t^��u��ر����A�����{G�
���!��wF���X[���:W�T��«;�2��Q�y8�G3�O�wb�~NGb��x}�ď��-+��rJ_��Щ�ʴK��w3���J�8U�Y_���ӖAvP�i�M���'x�5� ɫG��q}&���pѻ-�
I�AT�	�p	��L	"���!�I�t�҄��)�/,3�Y2E��ʹh�h��k�(#Ǣ��0A%d��,�����C� �hT>q����&Sbd�G�"�|�n1�!\�5�N�U+��ac�(c<�$[)<�~?X�UQ"��b3P��2<2M���+�7l)`z��fKN�h>��y��Zxi�N�X���b��]������W�#��y�clܕ���U≭3>'u�z�\&��Q:{����T}������U���@廝�M?d�b���b����!�Ew���z�[��|����A�� �KhN�����Q�����!߲��S�BT"u:a� ->[Ҹ%�+ՙP�:��5Ϲ��g���2y��Q����`2�����[f(�s/��K�����Y��bN /��˿W�ݟ�Z-���?�Q�{��6nߎ����24"k��@��d
s"7.��!bə�)HЀ|VV�A�BG�д*1�?���X���}����2�~�2��j�'�]���bQ�㋒�D��=�����>f>:���HՒ�n<�\��Gf!����<qT6��A��ɷ�)���1��9:���0�IK+3⒯����D��S����of��� M�~�vv�µO�k��Y�:V��� �Z�����]u���1� 7��-?/0�������R�����o kHVf��sx(7�X)�C����_L�w&N�u�`�������V� a�X�'k�.�|�$�e|�}��N��4�ɰ�~�*����Y+��J���)\?�2��9&:u��x������n�H���R��_#��S	�����U�O�)Cn�ߪ��<���*Z=�qrZ�r��M�����n7��F�e�A��;����9�|����ڸ-��0�HB��ͅ%[�� �N�^��m~j::6DX�6��%h60��E D���M��%$�d���!�Ku�#I�|��GP�����v��4�U;��w����pN���¾n�|zl�vJS�%6��}�
��˃lN������]@��C\�Ϻ�2N2�C"�ް��[����!&n:���_]�"V���7Y��K��� H�vr����}��$P
#�|���AP:���)��l-~YX���>��4���Rd�gU��Y�A~N��΁H�FW��Z8�kp^��Qi{�4�ұ�:�K�e��02(Akc���(�z8�:n��~W\�"��D�~�t���V�_@� �$�d��QB�/�0+̮io4�#� �q�ƾ��r��DP.�d��������,
�S%}��B'ҍ�['���2��c�=����\t*.�����4�d�vX�ck&��!V¹q��֚7��L��*{��u�iCM�1��N;�ΐ����*�>�SCŽ(F��􀩉�_���~�ᖼh����.�AH,<��`��*�FV�XH��LX��;��� uo�4�֚F�O/������=; M�NqG_Ц�:S�~���z΀��E_/N� l����KU8�ɲ���<�Y\rj�k����d1Ò%�q�x���9���֬�4�K4R@�,ա��8U����3O_�Tw7���e/%˓5Bo���N��d�Gb�=v\��@e8^UVP��D��{f2de����{��d1��/�,xӸ$^B�f���y�j�߿v�T.��2L����t����x]:�b��%�L��ڬЇ�^�����\:�Y�LKB�]��\y��E�G_\�(b?!^�2J[��<�+��:*E��w+G
�3�߸+����>d���6��ڵA
<�{�cN��//����y�"����b�HU������֋��p��[y����B�m|9���qc�x�z9��z��̃7���g ���ƺN��zr��J��n�b4<�M�7Ͷ��T��^h
�@�y����U�s�!�#���(6c�w	RP쮤Qő�Q��mM�&�Q6G�r�luY�� ��1��B�Q)����w��V�uU���v�-���W�7]�����ؓ�.�Ql�*��ƍ���e�#�Qȸ�Pv��"�J�_N4I-37��/-���1�$�H���f�8Շل�L%�/��w�@a������(��-gi>��);=Z���ǖ@�0�%,b�u�hk>j!���8�����7�� ����X�]���ւ�>Cm$��N�_fpV}�vg�T9Qs��o�&>M�r�|󉆺�$U�o��ah���~�`t�����AY�9a�U��� Ι�LJ�朮0�&n�\�q��@ X���2��%����n�u�v`���f����˷�J�ѻ�ԭA� Ӿ�V���/��"��-aq��b��O�ԑ��t�<<�v�d�hy>��W7vd߼����:��۲��p:	��8i& ��,o��n�db��a����4�@W*}a���0�s1]�*d|]	m;������]B�JwG���K�8
Y��2�		QW��Nk6ZXR���-&���km)Ք�9����)�iAAE�F�X�+q�7W^B�zRFh6��0ta^���#�8ˮ�烏���a��jT��[�`h�|'lv��c��?ʓ��>9�z ��.F	�6�v���D[�]v �.�&�[A�k�?�2��P0�ծ���iC��dh�Md=sX����ͺ@�FŅ��I��;��ED	���oʔ
E�@v%���K��]�@]�,�N�r����C��^fY�;qAݴ���*�x��KAZ�;�5�;e�6l��A=�ǛA��R��2~�_��ݡ���?Q=�x�*�W
@��(*���8.x"�p�8��aD
�Z!!�$l��F��wP�p%���<7@�� u�j��soy�Iyd�n��]$��Z����t�a�K� ���{�@_C�}����� ��/��
7w2��\l�x}y�\u���F SՔ,�j�s�c�*�;>Q�	���~����tA7� ��t`�J#���NwSɓ��Lu;�{H b�pU�Q AF?ܙ,�D��M���ְ*rF%ꙍ���!�Ͼ���0d��{BOG��?^JP�A��W�!�־��=�b��3P�{h�3�a�Ka�6�u�N^��� e�r�H|�0�/P�1�YYԮՌdL0��YY�m濕����B#��=i�[�8h�C�_��sSc�(yȦZW��w�u1-�����ދ&�J����9�;���b�:jz�f�b�)39�D�K h���������7Uk�;f&TIWс) TΠogg+��/me�ɪ��JIw�c�#?�`�UW��ha��Y<�
"^z<ȓg~���<|j�!�K�#¨���l��X@0;[��XO��Φ���fpD֡_�|����"���Ch�h[x��+2OJ������3��W�����gs�d�M�ٮ��o�����P�Tp�#~�Pź��P<TE#�\��`Gܞ���;���a�rɽy7zY��%��q��'A\*Qy�O��;�\�q5H�&<��~^��Y��Q�UD����D���JYa�{������m���}�kp��`� $�T����;����j�+'��'j���!I�v��|8q�J�`�zBQ���3�1:c�T�Sx	hR{�@-���ХA�����tε
ǭeB�2��<�Gb�X������g�pU����}nG�E?{����a4S�-��W�eK�~w���{�l��Rp��>ܭg�p[�2x~�G�d��<��2�Y�NǓ.!r�@���BU7�W&�H��4�!$�^7��f�J��X��z��M���ԅT��g�Ps=��č�m66w���j95R��N�*	�[C�Z:�K��5�RȠa���m����O)�&��h�^�h����Z��~+�� ��6۫�Sh�ޑލNW�L���oK���1&�@�X&��*������7\�� �D�S,��Kb3"�`���ی���X��ؖɤ�tT�PVK��J�7$?��q8��۸��x��h��Oa\^ ���Pԯ`�d�nsw ��˱nk!p0�IO��_�1b_��П�84�knXS�~&xd	��/������iAS��N{Cf8O��R�jٝ�'=X��Aڼⷒ@*~u�(D%����EJ�K醷��w�&�Ȏ�]
���lC�S\@,!�7G�J�,���1K��(�1Ǯ�"i�'��	OcY63��&��m�"�ͅ��6�j5�&'�f�G�kse�(��U?�x�Y2��������M!Y�EGH�2��xby�_;�-��#��?(�_�A�N� o������&�[�/V:��0`I��F����k�(;����.�jDK(CMR�R�?��p.`k�K��:��Q��\�
`�AcZ�oT_��ɬ�ɖ�ܗ��+*i�������Vޥ&U�B�.�7��s�0�R����;�3��(�U�Ә�C^�~K�t�"�z���~ulW���hv�Ֆd��K1g��e��g��i���@�T�c����5��8k?��#+Qg�ćumP�YԺv��t�R0�������K\Kv_ITto�.<��%�I�.CU��ZT5�*����ۤ$��`r���Ċ&%���=3p���,ѫ|3ss��+QZ� �ވ�7�gA�����!����ٱN�:`5%����f&����f�n>��SɎ�jg�O��5!R�2H���������������y�)5F� %u�E\'�ٍѰ���o����5����<y�s"�8�t�nʠ�h�=��D;��{Ry~�J,�LU����]���tO��J��T��t����YQ믓Ӂ���M
���ɲ���+��b�"�7��SE%z�9��I�[���p������/��H�J4'=�B�<����2�3c�*�bc���	D���$��:hM�˻��=�[��~�,H*p\>����g��)�(�̺y*g��T��PڳN��gYU�k>Q��۲�CR�R	��Y}y_��K+Nze�� ��}Ě>��;��z��pKYL7C��h���f|�b@�Je5nP�7.���9�X&��|9d����{�K�o��T�{��ۣ�M3v���ה/trs��LEv��� ���1`~�X|F��sWP�����>�{�YÇ�7���	}�H[�0��c ��l�;�[?"K���6�E���e-�3������9`���U7)����hr�w�V8A��s͙�|�^�"�(Tl��8H-�ZL),�q��u��N+�������Y�-�\��NP��~����y�I�D;��H|ZO' �f; ��{"�^�1������	��$o$|��B=QN�!R!IC���d������;��7�(��oo~f�룂��=?�?��ckB1�G"I�1G���<��^�Z�1�#9�Hu�\�/�ݩ��$U��D!�rmhte��~v]�JO��a5��{rlD��ɣt�]G�Wq�"E'7\z0)>��@��?"��1�T�Z7Μ�3�J�Q�;�,فy�2���z⍏�N	ݸ�I	���X�������~Q�m�,A�h-�3��ɘ\����ۯ]X��d�,�s�m��$��2bq��רU8�D��`ɜ�}��A�]Wg_7��?���e�s<e$��2F�I����n��]ܸ�u]\C�����d\�@����H��ϛ���o�V����ψ+)��Z�F�%��}J%����G������u���3Ѡ����]�=_�DrQ�gbd�<��
[��31�:�]l�;����j��LHA��ݏ�d��9�Pv-�ΗY#Y�����p�'��O�v@،UZ�f��іY����Q���&xQ����]��gu��A�Y�F��+�JQ`?�[�<���}�	�a@h5-�nM�F�J3�K���� ��T�/��k����F])9jiW��T�>�Dt�EeWT@zr�/���in|�i
Z���TB��ȭ�7Y-1�_btܿ���Zd%�K����p��r�4��nT�Äz��1,����t�
���Vp4�nA&\�J���2N���[�����N��$�X���S����M���n���nW7��[PeI[Jo~N�Z�_C���A��'��_��c�bQ�r�0pωc����������
0�ܯ��uȽ��S,�A�"�&]h�|=�.oZ����b�P`����_��pv�<�h͂(���R|����^����������T��3 ���K
鰳z_\JP�����h�1�_�9�)��D���^�e�p� ��=.�F���za�/uC8IJh�K�'�+�3�܋�Ir�J&ǐq���n	Τj�DA�g^߀�
txj�܇k�q�B]q&Y�DX(�J����_7͞_��gR�����T��^s[_��T��IW�!5�1a����;�WǵU*VԩmO�@S=�]9	bG�Tܟ"�RZEO����Xn���d���N �(-��9h@Փ����-�
{���
ڵ1�z'˯��BK,lN���7��]h-y�'5�j��5(��29>- �G5�rQ�Q�*�>f!�:�'�4�v�̓y���j_^Ճ�X"D	9�[����ZS��O�6Ȍ�뒰������z��#z������bҔ���5��~ZfIn0'�����F��3]��n�\pZqj�F�<9�S���g2�Y�,����T��
P��++��Ω�w�lt��ۅ0�v�]��ʬ݄��6��	��<��Q�� [�F�?��N��&
��?�)گ�`�Mz���r<Bv��"�#�e:�6̿H������<Ņ#<(���_���!��cD��A�;�R1RHO��(�A�1�2:����"fO��A{o%��Z\΍@�Բ���X�F�>KX_Ƚa�17T�5��>�"lҐ�C�8drJ�NoG�$�
Q~.��Ak�%��&��n��W���e�@H��پ�>�����b��������A"ss�7M�4O�������Υ��
A��-�j�4���hW|>ib�7�9�c<�R�ַ���ƌnKy�@���w�`$(|i7���!@/�%��>#챢�]��P `H���BU)6�q��M������RY���j(5�	���Fɲ_���� �^;���:r�S������w���r}XJ(�7FĖ"X�*��k_�;�u��Ҕ�F	9M��y
O��T�Q�Ku8��I麔����T��0�Ĭ��hL��N�ɉK��q[(1W��+E�0-��ޞ�3K)M�n褤�Y�� �jd�c�C2+@Xaɡamq�ި���7]�=1�\1��AR8(/ }+��\�Qx42'�|BEA�b���srstJ���ŜL�EK�
]�F'V�go�"т���'	U)k�4��*�<��
��#���2N��q����	�\��=��s��[Q��e���h}WW�_���%�!�/u}*j����u�}sA���΃�؝s{T��>�*��sp���h=$H�iZՁЌ�1�K�N���[���"�N��_�Y��Q>)�/���-;���e���qA�V��2��{�H��E�C�/V��f����O3�=4��N�	�D-d�W]���%��k��[�'�aSV�Ys(Fy�mёGq�+��H�}�O������~&:�|f5��@ǣ��2#_��KLh��@u�!�5X��(w5�w��#n+	��#��J������}�x���-�3�Hհ���o4�t�J�E�t�i��~hS��!�rݑ��0nA��-_%h�S��Z�ܴѼO���D�I�q�,�W����Vl8}!�g�>�e��2��{'������%m.�}8l��p��J�R��?����/8���7
��s|B����KH7%���Ttn|����) ^A�z:Bܭ�/��t�&Lg��n��byl�;��_Oʚ��p̌�ݻI��H����@3�_�<�
)HO>����j~��}MV?�e��)��\#EDAK�G�j#f@�Ơ�Z�|�px�pE��6�<�w�2�cpC��YL�I��u<e����c�ޞL}g���|��t�6G�k�\�aT;��e�"d}��~D5��N/���~ӵ�����2P�B佇�KIfG�]	/w3�����t�k� `�П*�P^n2�b����� &�)of��skxd���m�GݧCp��;V��]���t�~����]�ԝ��#|���8`Es���;RO������L�%�P���\�NgyLzΐ#���;��̚�l��qL|:��:�~�	�ْG�2������ࡪ����J̓!�*ܓ����ܕ��|]�= |\����7�^1xe�8�*j,
?n���N��o�&B����F��EƄ@e;�{������Ó.U���̵�2�oUr�nA�ե�0�ro'M?UL��	�X����6�h�~��p��]��+c�@m�	��V�H�,��^�eƩ#��lR8�u��lP���?�C��#���L� d;��s�����TԚ�-L/KU�A�ޱ{fF�xl�J2�m��ᦗ���_�/L5%�v[�Rj���}a�Ť� Xs��ɭ��T�#��h�?�����?ۤ�����^i�����*�xU4?�����*����uN�e���;���=Oe�!��8{{x��Zl:��:���7�h%���&_�,���mUpF��$����BD��f�}ȶ7��2�/pӂ�.ZĆGc��	ת8{�l�m�2�}�oC_e����|pp�١���ֶ������YSl�"Q���HPu�08�:].拭j�Յ�dd�0����C
�PTR4ŉ�,���OMe�1�m�V�����/��n��u���خ���r�o���d���/c��%��*��]}R�O5�<������i�n�xCh4h��OcT�f��H�F����S�o���"eT�>���2�� 1F�)�q�h�"y���%�٦i�y�}/�}��[���s0"�
�����0�x0�i(1���8���̽���'<D��7�vGe�����N�(�.+�*O�|�$)qd�$�D�.��?#�%읮�?�m���y�
��$0O�H�����@�@��$�5��dY�E����B�������,��|�����4B�Qa،�\��|9@�m�#	���%�z˻`�}���k���)��#Y���x]���9�|T��r�e�Ա��w��Ҹ/���<�f1%#���!=�۔R�Wd�~���i8:;�'�n5{+�����r�/�+Uiu�mb��W�o����=����_�x�`Y=K�-��%nu$F���Ql��(�?�����$/J�ywh���ƻ`����SDi��-R�3���]i:"�s����fCҒ�����B�GP��QUuS�ɭ�(�e�5��tZL#���(�%�L� �E-RH }1�[������ͫ�fq���K.37�35	�q�t�����	<���]/��,��9�1|]�.��ml7Iz[�̊�?�}P�sM��W��i�=f�ȴ�~g̪��p96� ��dH(�a�n�B�������A)����O|�G�\�zU"�[~0�$�� ���8���e 3X����v����=������&�vIt��Hf$�.Z1�Cρ���T:|B�:�J�s�Ϥ�k5S��cN��H���f_b�UJF'8U��z�;=P';���j�/¿+�S�c�쳡=, v`ʯ��e�B�qb�tHx���s�{���9,�`/��)��.�Ф �6�m�g�W��ʣ��]���+ҳ���C��n�S��g��2tm���P<�H�&kH�<�ﺅ��Z���j~�푭�408Ԍ�HJB;������u�Y:_EO7��|T�x~�Eؤ�9jZ����Trd�	��9�\tM$x�����!U��9	9-#J:�@�B:%�䁛���g�/:wfq�ZM�#�*�D��5������o3ݍS����vӻ(����]cv��t��mQ{��8�I9w��!KE��"Nɦa�J
�ԣ�Y��vM6�3c�MB���2�F��I�sE���勩\%������	bJY�d�\n��w$�P3˾�i�H��g?����=���\$�LZ��p�� ��ـ�`�-������R��h� <=�w.ڌ}{Mm!#�\�Q8SP�p�y��L���y�{��ȳ����Af�P��L���
a�"1��֐�'{�W �&�=A^���/��=���	����;��Ԕ�v:�V��E�'ޝ��&�,�Y�x�X��UO��"7-h�3�}HB�&�(z˿�U<��|�^�ֶi�э��+�Yp{�&d���l�8�E��1:δ�Y]f}�Ԥ���,����{ {I������I�I`'&�g
��!��1�.U��$�⪹�aS�,�f�|(\�N����&&��.�VF���O�ɖ!ݱ9q��I���� *���rһ���X��"gp�v�ȑ�� aV8��hA���o�̸�Z
wO���H�,`R��WA��S�
Xh���A�ZAV����_�h��֊�6�jݚf��ԉ���d����s�(��l>m�p�5F�-�����O���K ��O��c�=V6
�n���\��M�(�>3��� ���&�������L,�R�	�_$<���^�P��ֶ��SL���:�#��%C9�TfPh��v��{�U Q��h'Mb�ns�s�uC�
(-�}`nE�`q#h�e�C;N7,�
�߇��\5��5�#0k��ZX+iF;ӉŔl3�\en�7����j�+���-�+-�H~s'x!����E�P�қN�e��<X�.�|�]��ې�H�P#�P����q^�g?�6�L�bG$(rP$��!g�-�fH�ŭC����J�έ_%��Éx���0��R 7����)3�Ga(���	p�,�� �C�Pfw#�ɲ�1Y���[�,tg(xg�C���&G�ʢʓ� -T�̨6��x�)1�V\Xb�@����L	]rTD��sWp��ěa����q�DW���K����b����O�	��a ؍�Fi.���淇������>~& �c��`��Yz\W�`QhN��-�9�6C'�%��\� "?�_ �_q�A�F5�Q��2�S��F� L��* �52�ܸG�žσ��p�6E8RyT~:�����y
�����l� ȵm���ԄlJćM:����E~����5�^G;S�1�"�2I���X��
YH��v4"�mc�
�v�����r��+ߟ�K��9���v1��ע`� Ġ&�mC,nU�L�?NA��8�0�L�pڑR+��`��ڭ�Y���K�O�)h�@<�$ԧ"c(�EdJ�k����l�N�*�!������P����	z��!03�W�Lnc�Y�����5�s[�U���(�)IR�Y�j �w|\��Z<�e2�d>!"�J�I����=I���^�������Lr��R_X����9<ɑ�:Y�q�@������3�>����~{q�QM�Ѯ�7S�v��aAJ4}(�!�/�q ��G������WcA*���A'A�v��zt[�M��<�-E����Yxc�S�h�}j9��o�!�l����>��j(�џUE�

NA�&N��XJwÍh�n�f=�h�|hp�X�n�s3����tO�=R�L�	r�'���C�b��ؔ쉗�& ���)]�#��6�@c7�w����-n�3�;<G����(|��lo����]��6�5�I�M=}��X�y�#��sJ4�½D�/��ѓ�Y�k�o��"xU':�
b��j9�-J�������ݥ������d�Wu��С>r� �
�&�a��A�g1���r!�/s�:�2�gs|�d����᧸:��m����Sļ��/�kJ�rs��@�=��ړ)g�Mb��U����=���������Gp��\3#���>��&�yK�=g<G����}�)wl����0Y`A$,M�����6n�܃n��4����ղS�����b�1wY��݁���6�� v
�	8y!)Gb[>(5�1����ꉠ)�Kv����vu��M�,������w.��#��;�i��@.��ۂ��Wd�,) �I�ѷ^�a����5d�{�X=�T�TC3��'3\w����Lz.8U�К:���ƺ;_����e[��E+�H)��v���2��Q����a2ܙ�`���;�\uOT�Z��41�g�G��3�l�����oryii�8�
��������������-�u씔n�����E�5� R������N�3}CM�5|���+����݈�ehG��s$l�P��� .�eu�x��Gs�1`��39�c��.��W�㐽���X�}��-o�a,fZ��H�s.��f#��ʔ��֩|�� ���6��(D0A��K\������6��i3��.���m	=�i%A���<P�Y�Ȱɦ0�� `�YL���9+����
�2,ečN�X�8"l+��p]���B=�1����`z���ҷW������F����n%u_/\�)Μ�D�.|ff�'��g�9�Y�>ԅ���< �������7*hƢje�`���<�'��i��K�"�+������e�n��
�\0J����]$m3Ǟ�`�м�7ĳ�M[h���~}�1�����E�r���c�������Kp�r�'��y���r̎�÷��q��S�4[Q����� X�#��?`ѿ{�0{p�Q��X*vP�2��yL�T	�߮�%���W8 �М��>��7t����/++�ﵯ}
����B��M�!�Ŵ��e�;�5�̏�0�!4hc�5&0��P��T��".'@LƊw�g�.���ꦋ3�O%����d�	�9�J��@ڭ�:K��S���V���q�=��\�>?-��^H�����'J~��i�\1eGE�^_?.ً$�k�Q���ƶ��6��%�<�>�J��fY�q�!�a[�oZh�Ҋ�u��ή����Iû��Lp�*A���ݼ"#���[����+�d5���
5���q���T+Xc2@z7P��j��'��<�&)����~�l�1�o��]�ަ�)�#\�y&�&�n�e��v
O!2�&X�}l>��|W��$�U v����Ș��z���>Y@�یDq��ccTX�=�{��Zg��|�ƈt�����.��&|�c6����`l�VL�#� �\Xq
�-�j�t§9����&X��B=����(ys��Ξ���V�-���_���~��>���c&�2�� `"-��_ā�V�����	^9[%���uiN��`ޓ>�%��s�́ O'q�y�}v�Q5Oi�a	H���B:�~����9��hE�m�M�l'/�-�I3B���E b_A0��)0Vg���B@��)Ao" T�Y��5Jӱ��~N<Ğ�Y���d-!���p.�7�YsW)5�w��ÞޚyN(4TؑkʻW���('�Їt��¾�1i��O@u�2a$����GV�Z��
J3UŞt��,�	�%�>((քOӖ<����c(�4�u��P�pUC��R}i�l��l��eRF�̴R''��}v�B�ة���?f;�Ie:�$D%��\���i�F���dQ��HWh`t\��Z��ľ&~� '9�c�$���_�<�R'O�r�	�.9'�:�A���$<�<���ރ7��f������U���Y� ����ν���"R��y�}�)�~�/J_b��@5�\M �f��Y/�J��4�"�;F:�a�b�8�K/]�kq�*e��\����o;ʢ�Ni��|��f��d��l�)�ɂ=5������>AZ�1�ɠf�˔��8��H�a�{H�(�6ʈ��� h{� ��raUM%�7��a@��ŕ�<��}�q�	� �o$�H)�V>����lb�� &x#J��+��=�T[�]{g�`�]��	��O&e� ��E��?����k� ��J�S��?��i̊m.���G8sH����.�Ғ����塄�C��_�a�R�ѥ�%�@M�e>�9a!)H?WV슽����j8w�X4�v��e{X����
% h����1��22��*!o��5��8#�-*A�y�ɨ��谥�t�4P�N�;�z�<�C�QC(_���ر��P]�i��>L��.F��1�r�C�4K��tL)�߹S���`C����d&�?�p�yAD��u�t�.'2\z�^s��(��%�aףq�uR��\E�ۈm+u�jthо�o��0��uX���'/�O�y�X���F?��!��UU����C�#\_{�~�4�n�*O�ħXoǋ�ԸP ���#Ow�j+����,&"��G��Dҭ?[Y�=%09C���e���w��[[��	���>�Kt��B�'��ծ�\]֎I�t�D�B��O�w����_L�k�
E�W�aB`Y�N��
&bۅT�dn=L%�]f��YJ8����Ym�-:�̡�y���՝u֧��ǅ4�����!��`{)/����r{Lg�u��"����Kqs�GP'�.W�j������X�6�a�a�6��K�#%�M�b���3�	˄���ԃI�غ���S"T��l�|���w���D��B�m��U]8cW����5�ttgK���ְ���7M���R��#����q}�~�;��ߞ!<�T��ǳq��0|�l@.�Y;��;;E��!��H+C�렶�K�D�x�3�l'E�
�������E0W�-@�۴u\�m�}��t�F]�{���) ���7���b��P�3����i-빧+ѥ�5�ȝS�T$G#j�U� �sUo�"�׆$�M[:D�%s� BD���t��������@�͈'��,9��<ʜ4Q����:��5����ﯧ�L��0k1�˱g�Q�֗�-�s��믵>�y��9;LC�̐����O��DF��������E�f�)�c3������ ƺ�g�>\�Q�~�ǁ�T�h9K����S�?7��;+/�e_sD�*�M>S,B���=���_
�H���W��y��Q���]�պ0p�ǄW���8��w��D�t)����/,P^@�}�X}��B@H;}A����(6Nqҭ�v%�e���%�\h�i���L�ޙl�W��x�̭;߉'&�`\��Pa�>1��) )�Y�#�<��Fj*�	9������TBv%�����s�!�ALMg��M����ES�� ��@/�YKF͎�*��2�*2�wC��ת�o4��*��e� ����
 D ���
S��҃L"�4�]��eە����:�t�GƳ�C)��D���[G6��U���h�]�p�����9�\���n��_���8ڻ�tP~[tO"�Z���{��,��ȣ>o��Y�.��V9�X��0ջ�%7�풴�^��u�����e�@o%��SIcRtB!Lx,T���ͅ%t׍u
�b����[r�|���&Z���q�B��"�PZjHm�e!�ڼH� ���?2�#����2�_���m_!��CX��k�8����_��h`���r =���c6N��rn7���.��>�Ns����3F��rn�˅L�O	cHX�W�+�����	���ʦ��K�)�-j�N�����ꀚ8n�6������|�����t�����Hn0b���������>GE��[V�}"%�	�l�3xE,����
zyƲ˫��۠�f��d�^f�R毭�tRK��su/���=dE�Ns������UH�RB����9��&L�]إH-�Y�sk��4�HZ��±c��ˉ�z��-���.�\ĳ������;�����m��2��=U�<+��8����rw��+���t���J2�;����9V�^���g.(&[�g��Kȏ� 8�%b�ؑ[l�l��|� �7�&���+�L��$��J#_��.�Ls!�=�!����en�4��ڏ�5݇b��#����T�U�ehD�G�y�g
2�>�!�n��8=��c���1J\��cՠ���F�Ww���wӡ���nE8��8��?�в���
�yI��)"n�Uq��,������s��~�0M�0��c�|3t�H>�'�L���5����=�+eW�䟒;y;��P�Ӡ<Zޥ�oJ9���0C�� ����.Bzq|�5و���z.a (ŀ0��;Ӽ�l��Ö����=��W�f���u�)��oV��2r���I��>���xTo���>"�T)i�T��!���d�1A�z�U��F�;�(������%g(���.'��p�q�t$�i1��!���Ƴf$�V�&�,�[���c���v���US�[��[i�����z��d�-��X3Hy�<2�K&ck�ڪ��h�7<���6⡝�2�vW�,Y�{� ̤q~vAē��f'Fz�e��`�D�9.��ģ?,�[���v�ݼ��")iu����Z��! �14DF��f]� Am��CPƫ��-w=�q��6��K�\In��KBn��?���Ԛ�3T��%;����e�L�H2N! L�g�³������Ī�s>Se��-�G�@��Mad���I���7%g����%�� �I(�Ӫ �������@l�>�h~c
�,� o'MƐ9ˁ>ɪP��w0�ɸ���:ɼ�r��atC�����d< �[a����H*F�IVjFy\�|��*|�?���[���)Z5l�ԡ��EO�DS��l���=��%��C��0ω�r[����\hN��(5���W���}�O����o�*2p�P���-	
�2<"���IA3�����>m�~ǎ�ə��NPU�G��S"��fa�̱,�sSq�N��-L�k}���M�&i<��GU�Y�J�07����q6�J�o=Ɗ���6R"�������ZǍ�Y�-�@u2/�|�����]�ra�'��H����!;�D49%�t$cjfٛ�4�,!C�xߑ ���x�����j32��Û?�B8-yǯ��_�cӶ���: �b���N���F�s��
���0�R��T4-Nb�BP�L���wz_Z������R�})��\��Gv ��8;�r]{kÑ&uy�.�C�B�\�"��b����z�^S�()FkG:��/aӘ�]vׯ�lV|$��B���l����m���Y����>G#��K������J��6�@Sv,|v[�f���d��B�"�����1��)S�_�/����F[���x�xC%D��?�XYw��b�/;j��� �q�s�=*��nG��ʇxv��Ϗ�'ת�֌ �r�ȗPS�%�F�y����qn�@8'�ō@i��T�@��N�<��X�fH�^��T��[٩[@s���Q��l��7F\��ϋ���7J�X�G��7fv���--nl�f`c�Jv������/�;.�I �x��9w�}Vz���y#��݅za<�
ɡ�{֭�����V�*h��C�j!����B��r�2؆Q!��?��x�5����w�/��
�q��wd)v�#�}�v>�@Mb�td��k�f��p�H�H ~��$��"�q
�9#����P�	�g���T�x��t�1�bw����֖�?qh�\�0%^��ģ󗣚P,�3)������*$���f��
�ү�)x1��h(���б���lAdyC�0���j�XX�-��o9K��Y�M�No��4s"y����G_����@�A{m%�)[��8���w�%���-n�6��3B�8í��8��a͸�@I�z�\Y��8܎����$��c���!9�K�&e���[��Y&��J����yL}�Eru���
"�B��o�^
f��,e9�d�S5���q�?��[�ll_��Dنk�V�Z�l\�`�s�xlAT�C�&+fR��ָ�Ȥ�����;��^g�-��ݲ�6~���1�ͮ`�SsAˎ����J6��V���`�躞f�;W�v'�������
�Vϙ�Z�m�y�թF��f�e�R�	�#��a��Ja�;����2��Y�
Y	^�u�ݔ��Җ��z�]Y�����<��)���vuy ':Jw��3д���C�L�23�U&�����=���G�6)@��{��V^l`��kނgR6}ҭ<y�������j���4a��Kz�ŌU�	����:;��($��٪N��b��q��4b�]�E�9�w�y ߙ�:;�z�p��{�z��a��:v|$f׼����?����j���c�|$g�����Roh�7z��E�=U��)��F1"Nu�2�� �ʖ�f��:v;K+#V������y�M��7�6�m��jҭcWB�s�o,�`�R��-�.)	���\��5��#
If7"ʸ�]�"�[�!@�'��kC��=���]gNg�E7E��Y�
����������nOR�|w�S�{�by�Ug5X��@ȞBn�U���4婷IS��oӎlw�*(��-�H�M�����`�mtEU'�(�L\��z֏�
��_��g:��V�:�,cˡ!1�W�����]�}�w�K�����6�~g2M��|�ŞQkhh���Ш��/�(Y�R���2>H{&Ϟ1D��j�,4��M�p�챒]����F�+��
#o������O 2=M:�iC�&@Y7�v�D>������5v	}�V����n�\��xU��UH}j:XHϴ���P��-f�%�y��o��u�{��Z6e�\ L#�`��Ҹ�y^�/t4��"�T�li�@�G�yp���� "t�Q��#��M�!{&�(�7Q���u��_"B^�s�V��L�E�$�X,q�f.hG��������"�9a ��`�E�x�`�O1Dl�eA�����!`�������&�	�pFR���Wt�^�E�J��Ӿ�+�َi�j^��Jq�(�@�T+3�C�@�u�ߓ,���7,�ܷS��C�L/r�]���~�V��\�8�X��1",�:�E�p��|��L���K�����
'N�����o��٫Cp��
kܩ�hPPcd#�}�ں�2��d<���dW�S���Q^�u3����y$HKd��m���,�7��P�Fz��0]��$.Ý�o��+�(��X|y���	u��v�ڰ���:7�N$b԰�>L�Q�y�(]xUt&��yv5���ÇՉ�
��&��⭮�\���D�$�uj�֭�L9��ػ��ې8�$^���%C��x��Uլ�_y�aR3e�B&Z����+��ħ2GA�y�QoSײs�:�����u6M���T���Tݱ, R���J�J�/���h�.�VP`��yT~��IQa��s�F�^��k$�;�%���cA������Tcĭǚ��,^�N�3���ڣ�8�}������W��N��>L��'m��s�s�C�̷M��9���g`���g��,Gg�H!B��d�d���Po���ҡ�0ǪO�kY2m|eH9{�oɪ��u:�l�"F`)X�d8��%:�Ć0������Z�o����Q��}V�N�@�>l�m�_:��ЀQ$ZB���J��u��b������u6�gܝ>^�k�4����� ?�Vof)������J���?��ʆ�NQŝ���]6DJ]P�<�G֡���xLש�%{��Q\2����7�9�尤��Hs���N^�7*��F+�@rbt��ӹ����~Y�8t����� ^x>	1����j.�E4��T¢�TQ{��X����|}~@j,�rE�:�6��C�!�ea
"0��R�t�t��o��Pa�Ńk��A��m�W�q�1n�v����u7�7dTXv���7��	��l���"2�MA�,�;��֦�,�&�o�Db9�*_nր����AO��71VÕ����(��"�>���-�ȘR�1\y������!d��C��}���6]��3Z�5� �tŎS���p3�f�ki���&��|��_��f��:>�]�qfl�:�aܘɵI�J������ߊ0��r��B=.�WU�r�͠וQ:�m ��m���l�C`ICQ�LB����[D��J�D��/�z"�����c��`�V��Y$�A�X�� Q�s�4�(�p=��0s}��شr�АzY��W?��W��2$���s[�"����xͻhw3�K,l�#��(�L�|ӂ����r�{��펐�bZ}i�u"�?^��g��0�l^��������V�N�'Ł�,�M<B]Qn�黙uAZ�f�S��X���v��ի�ȵK�q���r���C2g�#3'���<?���B�(�J���+�6��K6����}�����h����i�R����B؆( 5s��.u����%����#����N�A��H4�No�f�&��yR8��ja�H�i��QխB������SpE
~��������D5/уz�W>;U��1w���I�6�<:hƖ�I�^{�����[id^����۰{Z�czg`p�t&�rɩ�a�L���ȶm"mK��f#�1�9���Ÿy�e8d7���G� Rj.���2����V^��{�FQ{�����Խ�+��Qapr
�6�4�a�����p�Pa#�����-� �9,݋�8.y��+]:���,�X;I�B6�V�����$��.����xj:��_Q�^ڿ,%��ЛX00�����˒BV��6ywffݛ�q�y�P� ��'���2�s3R/_��[c�8~�����{9��*
Yl�d	�y�˞(e���0��k�ؼ[�Z�8��#��S "�����~X5Vf?�J*�͋: �Z�/u�96t}�� �"X���x2Ț�/uZ���B��ʈ �޿?Oe�m��qݑ6-�Q7��J�Ԧ\_%^R{x!h��,*j!�.7��P,�i@��l=-2��<��D�E0�mG,-�9�
��d�/���d�I{V������ڷ���13e��:z��_yox)q��߼��?���غs�J��Pv��8f�ݻɶ[��A����k`��v��D`�=��VIn���DQ���!i�	}����Wg���ͷ@�_�k�6����Z��+��i�M��^ii�`�Y�`!)ť���5�[ۆ�B��ߩj��
���[U� Ypa��3]{�����Ǆ���P�Y�[�ҎR_T;�����(��Smy0Pc$��>�&9yEYT��~L�X��-�OҼ,��kU5yO���5�R��<��)�'P$3��|�_�x�s��=Ʊ�X�Y#o��it<Anu�n��l���+��+�-��@BRuҍ�`1��[zZ��6�MHp$|Uj�d��
U����=�E�ڑD jni��4���W���˝���_ݣp���Q��U-��l�qW���\-�*���(U�����
�D��?놺<v�$�)�E��L=��O�0&]�y[���^^�0x��sᚦ���p���{�EH{��o�����@2rǙ]��0���qS���&�򒔵]�90����r���f+V��e嫣N~Y��\P�Wi����.���`?�h+�V_W��w �`P�\3E����s�ҋm!WA�f!�����J��$@+���=V[�'| @Eעj�_6w�CHt�;�΍�T��F�ӌζo�~~x��TD�!���O]����1��64�\�a��w���%.���"D�	��>Jvx�!�H���p�f��C���v���Ӊ�;�s���Z.s15h�B~M�n�x<Ϫq�n˅��6-��n;�H�d���
���J����:>����®& $Z���+m%�s�al��|]��mJK�w�%�U�AP$��z1�@Vx��MN̰��)(�V�3��@Z��L�9xƴV�ӛ����D1��w��j���65
(�hB4����R�*?Τ�L���*�I�-�#��4�AU:��U��d�<w��^�.2o���|��+�w�Ұ��R�	VP�B��.LN�
�����_=8���>.�[��YA���8X�^��cU/�ګ ц�«T��l	#j�e��{����C�m�lύ���8�v�������ۈj�S �t�^�M�N�]S�l�2��3��"����3���$��X����|�Τ�v|�X]/C0^R����'k��f�Sf���� -r���)F)b��I��"��j�#���7�$��}���r3ׁ�b�-�4��V�b-D�q�1YU~�;���]?@1��s,K�֛���o��_KC� ���>`���u�d�����fA��w>�`���W�i�o��ɍ��0R~�Kჳ?�X��T&ǻ�[G�M|�.�l����O��Nm������~���?[\�9"eA���k��ΐpJsklݷoq���ъ�h'��'s���'f�	!ϯ�,��0A2�1�%7/`�4�~�Z����_C�yq̺f���{K�'��Oiw�}��%E�H҃�/a!��pD0��wR�%����,��b����Z���H���{���.�>�;&E)_ekYi7o�d��u(�1*,�9D����g��Y��(+��L�o9��?w�lE�p�rl����'Cg��O�y����t=30a3���И%�E+��)��k�k��oB�.39�u��Z{�ZW�۹�o~M�R�VS���x󲗽I^����xl��s�xh~�e�s����⽯��8�w��c���qUy&��7@d�� {�;�(�{��J��%�<3�Q�!H{�S�n7�w��>����.�
��?����dϡ���,!o�Q���������.��J����ʫJ7=�[h"�}ֺW 1\L��s�~�b@�"�� ��`�����j�J�Rɧn���X��3�裄,y
�/f�u��q��>ߗ0y�ӝ�e�9`s�	vO ���#_X�˪��p`,��etx�lF1��]��J=,|�%�������O��d?�x��Vu�7�Uu�٩��{� �8v�&h���$�)���F�]� L(��jGd����0��%�����]�Op���N�8�\�h��[>�[�p�!���]���'{�gbj�k��Oَno^���ۑ��gL��
7����tV�~)Kᝄ 6R\#l�i��朕�^)� o'�6�MR�rC{�}ՂL�g�Ug�抐�4��8F���|>NM��r�Q��o`ww����Q���y5��F}����N�Z?0#9佗1|��
��S�0|�w ��Ey�	wN6?�T� ����%�$t7��/ydm�ΤsOU�M�H��#�g(�d���|v����d�H8K��x�F썱K����чי`":��/wnT�W勘dM�+�_˘�5�@ʲ����`6��2�l����lLeNj�	��e��*�����֍���H��5�G"1=n�H*�n����[q�Ĩ��=��R���{"�疘��1�v�t�@���� n���BTǝ?�����8��_ʽۜ:�{���C�q
�hM�/8(8˞�J���F9��`b�e�#Pەdb\��܈lv
d�;@��V��O�[61NY���^Yʯ�L��/1l0�N j12(�Vm��O2����gbq���K�2ew$q}w$X�-v$'��!�R|�������(F��Z����JoZT�����N:~�4����� ���B%�Zɂa�t%qw�����RM�oj�:��X��aK��2��ߴ`���+8T��,��.8�B���e���93~-Bi�p�0�D?��	hX�C �V	��b�m"WU�����/4!�� �q�A�7��E�
��	0H�IQRו����\Z�:>�./b���?��p���C��z�������P�n5eG�y�EFu��цC�9ܠ��+{ba�K��2U�陛"I�/��3�x����3�2v��{̓�Ϊ�Ћ�� ��C�$P&�g��7QW�f���T�	�ei#��*j.ȃTۇ���0M���0�3@�]c/w�D�L�D%��+��; y��.EeN������"�=���e�Ń����N�W���U�=m��w�q� �H*#�c�	Xbk����D��Dl��ҵ}�1��Y��lL�MԸ#�R/o�Q�M>��R�E�j�8Y�f��x��ڼc_�f�<9u��jW:���/U�ݟj�E���;V���I�>� s��r��0}�O!т\MaD`Q��Bt1k������6�'�O�B����n�pB�l�����J>��L�s,���T$[h���V�j�-�����EE�� ��%�eځ�.}h6����&A1z' ~�F[Hd�:��7u��)U5��i&ɮ�*#~wG� ��Z���i~��-5���r�{O)R�Ƒ?�����G�@��Es���UǟD/����Xsڔ92'Yq�s��\����Ea�����KA�'q$�ߩ�k��TM+?7�"�v8�kȱ�����RPV%޵ǅ�.x�M��_��bƤ!�����K�辦���5%����!E��$`��/m��;�$�~��~;7���(S�%���z����S�����H+*�<�/�9\$��r��`m�b���
L�(rC�u�c�Ci+��-Qq��b�؅!�p-�&G�if����$"�TH:DO�4���pcV��k�����K��$x��yN�[���+(�K��N���h��rsE�����=3A�	�m���@K���� j���/���"���"���b��Fқ�}H���6BW��fψɝG˒�2
@� �3����zX���p$Tk�&��	��
�X���`�7�E��Ҩ|;/���,�`.�Z[O2��_�w2N��PC��h�561������::[#��Js�[�'⼻���UXi��{#b�/r�����?�L'���̓v���7�O0;k�4���X ��󚄫�_��R�Z4f��=�Q)��g����9&~��j���3��`�E�c�����+&hMY��WP��ɜY��!m�LSi�(�
����?��4�~uc������n����c�p���˙u��;�
7�n��M��t���N�e�Y��ջ��WtF�"��^�В�L"x��H���h�s4�he|�&V�qwfc��ѱ�d���w?��W��o����� ���Oo�h8x� /N�B!$�KG��2�P��i��g�m��ۋ������k$4On�����*��6��Y?��$r�8H��;��(�a�4�
RÚ-�� y_~^��JG�h:7}����BL�E�%�v�-o�q�h�U�5�0�M����R)���1E`mЗ[����F�*���|ww�Y$��u�H��9���K��5��%f��L�˙��k����L��V����|a��8��B�$c�]��r���r���4��YH�����#t��]iC��߰��#V�,r��b�W����.W��;��Ϻ����י@Ŧ����7�X��:�`#����}Bw���ֻ���N���9�ߋA�:�ܾ���\B;������sP�pK��b��~�XE�<{�p�����A� =����Z3�p_��X�Y���|���d�l�2�?�<*���A���#!�+�\a�eUqi÷���/Ya���{j{�K n#�����x��;��7�*|y�����3|�Ž`��*�G��?�)��UpT��3����C.*W��t�"$�S{�j?ZTA�S<nAOb MN���ˎH�aP��#2P��'�ϒ?�Z��Ne_�re;Ah�)ލ:p�7�d�zo0ד��'�N����cm����Q�A�����9<Ԣ�Z &�����g�aTzQ�_ �m-��mR�Ɛp��s').�O=�M��o�',���vh�Z�{�n}ݙ��9�l��2 �	M/ \^��u�YJ��곯�{Xt�<u�յx�氬KC��ojDc�Q���(v��:}�RK�� V"P���۽׺�Z���!}_����򭥜��Q?X��1��(^;EtY�g=#�����!H���� LW�Z�P�~��G^�@���!�ʘ28t&���J�F�)�.�:��(��4�kNco����S��U:�#��v�Eאw�K(�|̚�-��'e��<Z{Fۓ�uq�z�~�\"�b��%��n��s�Ԡq6��X? �����R�_@��ȎH�P��[]{[���:��̓v�+w����v��9X"������-�N�|�Q�:K9���d{�R*nu�;u��nG��֗�Z�?%ޖ��w�+H��v�3fl׫�<���*dAXL���U�\l��]lďu��-Ō�/������8��BcG�O��lx~[��]UJ�[�ʞ/T�P,�C�q:��u��-s��O���{s�lRa��:3ȯ���+LL�����[Bv�V��6�x̒,�U,������ܱ3	�����+%tVy_u�49L��o(�;�!�a�,@@[b4O�)�

ה��BA�L�<}��ʧ�	Q){��?���0�)jla��%x�v���3��O�0:�r<�O��x�^��u_�^�t2N�4��C��)�Pi��oY���W����ɹ���G(�U��3�G �ଝc�zh�Rɹ�#@D���H��gXY�T�L�U^P�jx�B -��j�-�Pb���)�挎ds\��&Ń*�d�2n�8&�6�O ?�#��C����e�1wM|IX�'"����D����+n�z�]�]:X@�T�����G�ˬ�,)��N�Ç�گ�G?�J�0����	��ަ���b������]���(��U��2�Ν̹Bk�N���!��8δ��@�i�7˕2PV�3[xv�#�D�{0��J��N�Xj3���U���:���3�6pA��:��4���s �q��B��/�E�P	;O��i�@��S���#�����J���������HTp�8$p�F�;���A$�k=��q�VQQ�&�9�WP�G17FQ���I�)@�ža�Ч�|���M� }���O��l��--��ؖ��us�����>Be�����Ȧh-�>�F���L��}�?S@IMwJ���J;�!/M��b�g���dإ�:�Q�D��ru���v��oJ��8V��`i$�`P�x4.0��"Z�d}4G
�ވ�U1���`��0vB�hB�'����"�sCW�����L����a�'�[�q�E��i��'� ��g.n1�>ݜ8��>�z�~Q�LWl��_�����"��N���!�����y����b2Bp)���(�W<���&�$��i�>�T�0
��"��$3g8��	U���	0� 5ڸ�~2&��b&�t�t��6\,��� ̐15�*.�j�-���rv�v��3��� ��v�V�"X ٵ]�����1ZKp���&^�iq�1T=�N��4�j��rx|H1,Z�}�=��N�����M׻�8���a�v)�w*���1&���~e^m#�P�_����n��.0�o�G�X���`���i�ih�c�bGc9A����ktNѨ{мS�x�`�L�R*|�]��G{y�r���9�,rK�S�p�!7��6K���r|b@F��4?6���T�WK�Ӵ�k�gE�;�6�7g! �9�J�d�v�R>iN��4$eL�L�3�G�	��13�?�Z>�ȸ�xT*g�5���D����W[�ky��{B�������)�^ܪ����Z�]�Ű�m��RJ�(��S={S���pXy�?�"����קF�Sr�&D��W�>�`v&�	.GS h��)$���>>���+��%"�`�Z-����0Hu�2MSG���A�y��*�,�����Z���du:41�)Oh�]b���i��.��ˌ�4����P�A;��# K�}��
�N�
�\oAZ��%��k��g^!kV���Y>ˍ���%e�A�Վ
2>�Ԇvȡv��)��/�E/PH�`����Nac��$�S��8�c�|�I�	�4o�ZC��zsu��1��	q������ؒ�C�^o�U�ً�.�.����pr�n������9og�S����HҊ��+��:Y �����Y��"��� <
Hm*���nV-��D刡r.�(���0n7S�I4��
cԧ�T�G/���� �<�l�J?�a�[	�ջ.�u}��b.� �虲�{o��3m���&{2��8)���7�Z������|�|3Ӳ�{p����CV�כo��8<ִ��`!T�?<|D�W!pk��y�(!��*��"�W5�7�e�u�H����ϟ�-��=��j���V����Gch�PN2��|�A��GrSq.G��qя����8�҉c��ĶG�������$V���I�*�GMֳW��/��۳���O�ٔ�I�·yїr�T{4�!;����C~Ԫ�!��!-ԛ=]ޏ�$�&:��ڦ+�!#�������s�� ��$7M�J��d�5������vD2J��Eᯬ�]2�P+5�����$�edI���F�6q�d�D�a
���w�Ă����G̕9��n�BDe�G�-�A���j��⻂����vA���~����m����DW�>A�^H�if��u�������F!T0�Ӏ���,75�IdK��]6.���̓~�������=�}�s��I!�yy��D�n�!�#k;s�KUX���H �������5��ˈ�E�w���]�iW0F`\���M6�S�(�~S#s�g��|n�s��d�8���2���-2�T��*y�-�ӟ�KE]M)n�	�h�{�|�)��p~�A8��ׅ���!,�nc�~��t=#�'k4ק'����j���"/�l��M�ȕ��?���<Fa�A�rH}'�{��aBšv��u���|H~NJ��I�P�گT�d*��v����l���s��R�j�Χ���{^p����"B������0�A W)�c��w8�ǽ�.��l��6
���9ւ(�����j� ���9'�IYㇺM��h#��<��������g�1�8.:wR/tG��Y)Vg��!J �h�#���[��zN�<cB��A�Շ�b��\��}�O�+t�E&ttZc�'r/.���w`����l�{��\x?�6�xͮX?t�0�W"��8Dm(ݞ�^yM��m��%�?&9�3��ms��?;�!o�>���ydv���������5���=n�q�KN�烹�AM*I��z>��_ �6��	c��+�l���^i9<��6�7�Ee���6w�*�4��|4[r�R�v0/�$`~"f�Yk�'������3Y��T�$�*�VJo*���	����EPL[�3��� ��@>`H�U:3���L��x�w�Kז{B��d�(t�����K	n�󒺩U��8�z_�I���z8g��k�bKd	�Ȋ��w뗿w�W��ݨ�X7���@��Gd�.�A}|�_b����b�Y�Cl�N��<>�&R1��%>ee~���g��$e�,nR���+Q�<�2�{���ࡲ->�F�Սo4��<��;<����H3���a�
]o��YsiM��߲]Ө�Խt��EUPg:�t��Mg��Q��	�O�I{g�f� � ���M���l[������(����rǶ�c�g|Xi�Ǘ�O-�g��=�z���=���O�w��R�����_1-K�ȒvdZ�ODj�p��Ռ�!�pV�X��'�\�۹��'�?���yfŘ��Kģ̍��U��a��E�
�����k����[݈����b���P�F�lE�ō	���m��&��,Z�r m��b� T�K� �ɮ	���ɫ%Lj��=�o�R��P�8�����+����ŉ[2��L���(<���������(3'*԰��m���+=P�
���
�[71��xp,���k�a�"��"+�B�ʮ����=�,�f
��YU��������ŏ,��iz�v���W�0�M���%�Q˽�^�
+`��}�����(4�fDwb�+Pg�DBz�y�:��u�J��RDe��A�3�Ny�I�J��J�'��N��]_,1�׾�A�y^Y`����U<n]䃔�%U���auna��g�V�'&��}f2����9"(r`�3���f��J���w�W6�o�L����; ����P,�.(L���1ŕ��!�W�l<b꿇�������p�&�Ô���ͧ9J�#^�J�Q��������7kר�� �=��>Z�xi��{��b�u��m�&Z�����<�_	A�m{.hx�{<J�5u� �v̱�mK�0���͓ջ�p�SHZH`�����p��Ω�(x���;�\o��!��+Z7lA�[���OZ_F��ĸ[�b��3�Xư|�l�t�� RJ!!_T�`\E�q
����[&���i��R�=��P�56W6����ڣ.�ix� 0�dq��h��qݚh��(zZ��%(e	:��x��[���h�`�6ǔѱ�<ǜ���/���A}�Uib��LE}Ta^+ꏋ��J�f��HSrV���oM�66=n����7!#3jyJ5]�!\i�������*X���Ѧ,�̫3��0�r׏����S��{ȴ�8'�|D�Oz�9X�rn@Y�)��5�KzEM�����rDlj:J�4�G�=n�(0�v�g�`��Q�O&�w�bo�m���m�5��Z�8>HG]�)��_��ģr�o"����O5�����=������u��rl.� �� .��I�F��O̥fݪ~'S|k_���8��6K����cmT���P��s���1��r�9��ϕwG��tm"}�q��˖s=h�]�&��~��rhnI���%������6XD��{��Σ+ �h�A��N�q�@ �ZI��9����tו�q8W=��10�������w�m����Nsf�C��{��Ƹ��>DӑDm�m�3���é��|R=�����?�K��X�H� �{�qn<�Ei���o�!��u�#��hk�}��>PyA
�����f� ����L�����xW%�M.�Ê�֤��2��Ji���   ����M�n����q,�ʄ9�Y�c��ܙ|q
�i!��i~�u9�F���^"_0�
�R�1���>.�7����1�P\PL�Q��It�Y{�������&�/y���"]��e���N9�|�»����[u@�/Փ]�"N{���NLN�0�^�0Q��,��Bl�N��b��V1,�ݧA8V��<C���4�0���+=��H��7䶄I�cI��fv�d�����{%lc�1�C�pF���h�׈j�rx����~0��uJ�[\}�=�b�I ��(	�
X�=q��Z;���z�ϓKP�9k-ƌ���B�Hp�p�!�e+���ܿ���|�ʇ��D��<ie�<��ύ+���������0+C�l!4 W����2\* $�Ũ�ЇdZ	���o�ٳz�⚋*6��_N륇�}c��[���0�qEQ�1�!z�vb�w�����k�Ck�g�d\ݖ��!�~]
������k��à�A�1��/�ȋ���#�U��1�|s�� ����ځ����h(&���+r�qi�����|�;�O�ՇdʜtZ���,k��b�DʆC
�k��3O��\zFKH޷X:_I��<�X���G�5å��we� �2G�&��JrY g�o��]������pL�J+�W�l����]U[Ꮘ�9l֚M�P�A)c�K���O1��<N�à<hl���Ծջ[�6��K�d� ����-�$*�+�������o��25�/^ע>���2��zOZ��h,
�Q^�v�R��xd�����sD�}=��'VB^� ك�$�V���}�$zƹ=>d�5Y���!��F��mr$ö�yƏ������}�T�[W���]�B$�M�𩈸u3d[	���fO�ߗ�P7��D�w.'�^&a����zέz�����?ȕԢ��2*מg�2�y3pԹ��i���n���r����q�@�v��YO�v��!���Qg��Qh������5?�>�����g�.��Fy����؊a=��j7��c������`aT۝\	�s"h�3c�|�'�)�i���A)�@t�3Zx�Tn��������dC�G㩽B���B���3݁l|�?r�+�aZX:_��Ǟ���[��������
����G�13ѾS�~��t�PI�a�i��f�����"���Fn�EMPHx��:�v�#t�u;:�K
�8�S��{l�U�s8�֩�-���3 ��վ��t��D>���4.�{���n'�?"xd��-��l?V7
R��0
K�p��{`/�*ieJb5�^��������_��`^��q�=iVA(��z��,VQ��
��<I���[wz� ��ۚ�]�Rn��}�t'��_(���'�d�m��fo��-���Д��O'>d!�Ԡ��5y~�-m��o����!�4�}ڒ��}޶�L�s#dk�OeQQ��8�r��E�%��!�3V�[S�U5���j��S}��|��j*�¥�)��j&����E��W���ߘY�^"�����};o�~V���s##bٓsj���hE��7�Δ���ʯNV�$���q��)���жK>ASY�� ��|�n�y��
}|?�1�H�b�p�<~ 7&ߕ�F�S�?���z`�^�f��f��%����o��`�^�*�֍T)([K�i0E�,-��P���'r�OP}���p�3�dwJb��D�v���2-��.	
��q�7j�g�%�����\m��T�|��z8˱9C�/�(1&|.|��yw�|�`~o(����Wt.���&tޣv�TS��m�X�Y�	���7���������|���������#̲����3��L.�N��Ft� "ё���/��5P��+�78�۾��c�B	J*s�CbFM�_Ov�WRs��޿�(�{5�^�=�AS�\
jL�.�����W�f��|G��S"�1NEZ{�~/G9o��6��O�DG��d^�Gb�f.N$)����~ҔV|���`�$,�g}�>�T
:��16D�"_����A�T�-uC雄`V��h��$��/ڄ�z�h��0�L��!�lлP���`.q��IO��Q<gF�N\{�A^�����oh���ċ��k+P�{{�C R�o�gW�Ιr�g%���H*���/3�_�6���t�Xɉ���
d�D�\��|tS�ƴ�&$��E_�΄L%��[Hn���؀+�I_x��bڝ��������i�+a�r=ݞ$ʊI\ ��\�����u�J����~(�tR�Q��p�Sk� ��4��;ѓNB�iWy�V�K\��~)g�;W�utέY�k�/Σ�Nv�9�� ��P�6ʖW�uJg��P����S��4AKw����N�Oo'�t������R��&b����(��H">�i62�F��Ǻm��5�B?��v�NU������6�5��(�f3Cށ��T{@. E�&�ώ�6�U@E3��v<;y}b���}���:U�_��|2'�n�9��c�הp�?]a�J�+��NM�<��fH'ʶ� J�	�ҥ��ـ��ɗY5��ؘ�e��dq��`ތce��0�'�X=r��m8`f��E�4e0X�Y4
ƺU��̭q�6�%�/�]�.��> K^'�,o �0��Q�ڱ���u[����L��hiK�sd�K�v#慣��3��d��5�}R�1�	P�eEW�)e�)z�0�R����_�<�_��KR��ۘ��i:�͎S��\�����k��ȸ�8�|���ߜ�%��Ђ��!�:��*�mU���oZ�+i n�WBÊe����G2k�� ���k$���W�m���*�Ћ,�V		��gZ.$^��*��cqh��B�!�ݞ�|p��0�(,C���ߜuT�BH��&!ly��q�OCGt�1W����(�ɝ׶�)=~��E�4�;B[Qz.⠞���]X���p3t�%�2X ]nfĘy"�<�+sZ3���''�Me�GГĲ��7b��0�Ҿ�q��m��"��Dt����B4SP�{�pbo��s��׸�.��	�����{��Q!m	��ݛ�հU4/;^���)����Cb=�F�}L�PJ��ܷ\�'�6�&�ֱ:�`�گ���k�h�+��Qu�&"�ـ��	0?�C�yQ�z�d-���%ڏ�c浭{��=��zm���rKQ�'�h��7�YMD8�\�꿏�� �m�Dc-,�p+X�垢�"�;����~��X��}]���p�x���`�99	��9� o�GE� _V�vs#��_�zd˝�q�� 5�~�YFg�᱇�P�,7��N�y��L�!~� �ha�2��/�K�'ڣ�PP)�2L�08I�{`�+t�.2�+���c�互|�N�����bӋ��ɶ~��9���
M$,�nm'/ړ%���f�'$�fЇ��M�Q�<��oY1`���S�L�*#�Z(X����lJ��]�}3���J��'�,�+���������ڄ����X��S�W�S��U�4��aZ<��rW�n8�L�K��@Y=U�j�]��-#�?�|O�\��_�Z��eC�,4Y]���)��F;��s�P�Aޢ<�`o�����.���g�O�T����`��V�=���==zS�u�����Nw�E7݁�V�G	�)��NJ濋�V�j� ��
�B@�3�����V���NƟ��S�*�oc�Q8��Ǝ1bv(���,�i}1�r�2�(\dF��o�E"?�C]j9�C<ԚI���4'A# �J��-?�����F@?��S�`5�9�g�z��{|�����}F%�eo:W�����@��{2zJU �������K����@L�e���z���{a�`�y�� ���b� �m1�5��`�b��� �1�
�[��w�Jjib�o��`�T�d^�����Iv�`�l�C��>��6_N=#�2"��i3�7��2&���ԔC��je�R�Nt�9T^=^-�KuH2ͪ��� �F� �f�T���=Q�]���&�G���5�Y�X7���Z6�@nf��"��^Gx�n,��д��gs�e��N00O�v�@��;��Vt_�ӧ�Y���~�m�O��ƓT���@��F-֣�~�7`+��+��89�=�ڼ���?I3�*����vo ����%��a��P��Z��t�!2{���v�K`(�	U�~9���k��"k͢���=�� I8��{�E͌��fe�V�¿��ߐ����|[8	��>�o��vr���ӗ���P�iͳ����u`�2�ma����g5���À?P�	l'
B�ש�ڙ<*� �������?**)�[�F��8���
���w�(��0ÒQ��_olx���O�̸��z�B��57YwVh� r�����k9���W=�IZ�[�ۘ�UL���@@ک������s�Z��Y0�Z&��v\_�a���6F�SAҸ�#�I\r��Z��=
�`tn�*�	�D�6��Yl;��y��)����ᵱo����W�7���*���ԓ?l��mh����M�.S6�(S8C8�O�v��'ؚ3��$���z ��C�_�c2na�ͽ�L�TS��/�Ƚɮճ�7�g�Άn��C~H�b|�7��Ӝ�)}RjU��Ě:�{��H	B&�$���(�t���Y� ���Nz˨�����n\�.'d����5nC�2.��}��ڽ� ۶���N�p-�;���e�U5u*`١2[t��L����]p�ד)�����T�I�`v�c�)iE,��jIB���/�o<�^���P�"���ʮ�#G`T�]!�85���uh��B����<��0K@�����G��ll�x��*�c��yP �5�PNV�p���`�*y3 z2}�GCy���"y���/� �(���(^?1�~5�?)����N����2q6�ԉ�M �L3�.N��]��
|q
`��tנ�����)�G�� m��@�@"?`���h�j���OB	��Þ��]�Y�5���8Ē�uaW4�#����sh��uz�Of8�s���9�P]7��P�y� ��lXԉ֤iш3�n4�a\҂:Y3��
�`�@�&��/lR����]�@�)���9��pE���Y0�oe��`RD�r�~Y��{yVv?!����h�Z����ac�U���j.*L�	�-�>j\H��2��a)h;D����iwD�YR�l�a&�ڋ��j�Ȭ����Ľӎ��]lk�~I+�9����4�S�H�go"w�r�b#�@�`֊ds�)(>h�z���NFnP#��H���^!�[��/6����"i���e�!�/5�嶗'[�H��uK(��/9�9ˁOk��`.�n�n"�<�ݿ�-}u�io�77���x�e��] �� f����D���O�vˈU@��.�C���i�� nyC�h��mg���r������d �S�o���V@�c ��ؽ��\��(�7qA�=i@�f�l��,O�;os�>ʕ%��7]�Ɛ�g�~t���Ƹ�z���$�(�eI̸P�4rZ>%�(	�"��,��.�$�NN ffӺ{���/Q�O\���K���ë��`.�k��VAR2b���ª��%U��ku�P��G���P���?��f1h����|_�ش t��y�?p����|6�;��a4��z����?��_.a�ͤz��d�Qa���ށ���)���:�-�Q�]aŘ �9�:������S�Ӯ�T(���zKRDC�8;o!,�����!�D�<��̬��G�[�_w�ʻ�A~���2i
^�dx6����Y[����̔���7����o�Ш��Nw� O�/T��b��a^�G)F�6��9&L@���^��Od������<N���'��V�ÞF�┷9D����O��?ux ���_�W�ul������-��B��'�r��X�i.��w�7a�\�Fq�&�GN���D�nݾ]�8� H�^JG��tMj�܏;565 X��d=���޽�f��
�MUD,'{؀�������<t��NN�8��4"6�,S�� @Ѥ��E�¾=*K�*$M8f��e���6!�-¿�)�-Ъ(u�YD::��(a��V�hE�1���wB�Y?�e|���H\�l�0g	3�Gy�z5���Zύ�0I�L��d�/R����qd��{��Es����NVy!(qa�-�R�{��U�oX��.Yq(�-����J����:�x�b�l�z��lS%uJ�(���щ�~���p-C@���]����ζ��b�m��/���Y��v�U��}�g��_gK$�P}u�V|�"�jdRZt6zt	�Tq��7.O��˧nT�7�@�;�f72���⛎�Z G�Kuȑ�ey���6t]�0��5�!G���8$�q֟�Op\S��Ow{w����2�<�b:���x+,����������c�g\����%h<�*�6X#+\�C�%J�����t�#d�����,�,�
lp��!na[)de`��\�l��gi��F,��z8��gi�A7x���cB��m�Ho�5R8��G��p*��w��	���&�V|����,gjĳ��6��[������uI
'%ת���_�k�L���2�m�[qԋj��x�<3st��{�"e@u���s��|%LB}W��@3���Lر�yt�;���b�R��+V���׮4��� kYK���3�EP� ���(���SӅ#����My�3�z`QTT����H�<��w��Tȓ����R�R��[��!��6��T�W~���喦|RȪ"�i�"�q�D�nN��bN.B^6p���e>�j�Ċc���3Tpe_
 �$0�Ȉ̙��2�{�sd�ȔbN�Y�'�����G.4н��Fs���N5�w�0�dW���t�&ȃ�f8cąD��x�_:C~�p��IZզ�pM������Vwd�_�cA��g]d�m=|�O`e6��:�To���Hz߄�p�O*3 9� ��}����_ppv^�pīF����2���b�J�آ?�<�*2�})\�ʐП��3֯�!ܵ��W��1E��y;@x�k��-�\HW!Lw�cl�}������E�p��u����E	T�C��cB�ݮ��� �0p�EP��3�L�)Ig?�+���nń_͇�/�
(��4X�h�L�ܱ<�(Y6d���"gT6�m��My��2f�E���Y��*s��#�	�lw��-�_Mg��91�����B���žW����a*��	�O��"�ʹ]��O~���s���޶�y�`$td/=��A�R%�n��"Z�K�z3/[x�@V�C$V�PK����� :�,�z�����¢8w����Y�=~a5k���m�}�Qᾚ����S���Q'�>eS�0X瞘�������g$�p�7#ǯu�؞�>�����?�~��m����~����[�M�ut[(�Q��T�E�>����[#�T�f��M�t<eC.����;ۉ�d�ڼ4]�%�jn���g��2;����Ęd�c����Ή���<Z�����dx�Y� V�1>V�P�X�4�E�%���w�U���z��o��+DW�{bײ��u���0�jC��;ҽ3�MG�B�ч����:�;�P�bl��t_��qۂm)�&��W/0[~�d��
Zj����Z!��ğ�=hy?�����(e2��'$�#o�T40S�g����d�f�A�(�W�O0�q��Q�[���Q�`	6�O4f�� ~+e��Mo��K���-� �D3@/<(}���ՂC�4�����0OS��DA�TzA�*���+W�\ID�1���i�s�p�rbu+����C��Rc���*C�~����a��M���g� ��� ��9>���2����2�@��8Př_EC��:/�u�b,���"�� �W�#�*��-�Uj�3�U\�"��A�sJ$�(�r[�u*��[�k�%`BA�,|�#���
�Z"Zx�x)�t��I�*�.���p���L�J�{�O�Q�%�6���$�qC��l_:�^��2����^0r.������CWs������n��:--�F��MS�a�ޚ�65�g�3�;Æ�-0�Rn{��q���'\3>.0�`5�$-��)cD�O�gx1(T"�Ӑ��	��֋�ɑ�*�빌���3I��(�1^u�i����󕙬Y8=.gR2��2�gBCtX����5�@�)I N[�����v�k���G2���~b�d~�Hg���	
9:��J�ـ���;�T="��s5O:S6�S�<<?����B��8g��Y�M�Q�V��Eb�	���3�A��â�j�K�;��V�;�6�}�&Ԁ͆a�w@��o���!��~p��^�P�%�W2T���Ycf�iкm�����K�����"ň��K�����Yn��.���(�W�f��gȮKG��R��s�"KRm�k�،�~���
��M�/���&u�>x�u�M
#��-,��D��Tn蛯�f8�����D,v4�;�U,�s��e�Z��l~tn���(��`�I���),�����kS\AsLG����Y)]"�q�R��깓�� H:����������ݳ��z:
TL@*�3G��iϋ��=ʽ�~I*������(q��&Ȧo�K��R�3��Gc�ģ�g�0���}�1�1>����g���fTUˮZ����k�n��$/s@B�[=i I<�9�6��>Zv�k����]�·�ahn`9؛��[K]e�F�qCe0|�f���fĎߚÓ�-��O��s��`��ϒ�ײOv�C��WH~�,�ST$�G���(�w�ua�sn#a�V}}��"8k�pG�B�@(l���`�G�0�EƹAM�Ts�}���8��uBg`�\�(��*
��C����k�E����Ό�yTI�{� xn)�]���'��8�ꆏ؍��6��ָ�W%�Γ?�hQ�#Zvoy��[2SL���]��f\��:X)���/�4C��9��'��?:�x��V���c�s�#�f������ξá�?�F.���K��ҡ�4А2	�D�,��	�<uZ�8r�8�H��|�)g�x��y�C�Z+�v�����5l����)�-�4A�W�`�%*��i&�T��lp��t�Z��0�j�ͽ�>��.�Ɗ�W!
�l������H�b����������b���TE��зO+���[�S�W�SU�c�/~�P��o�[\�I����2�b���׷[��I�ׅj-�*S-��V,>��W�Y���ȓw0tLW.�*��3՗P�m�S��U�Nd� g,�@� k1����(���,n���At�����2��	�ۇˋFj8hG�!&[�}U����E*�)��ջ��ɻ���^k͔�Ȟ��I���z��.-���r:��U:�粍S#�?"у-�����tZ�����]��w�����鞢r�����0tl]�e|%�}T�� �2�en����	x0F� �:��<H��7,���vO���
!8jANr򹍈y��zk�Mj�`�:'���yG�,(�QLE����.�gS��;K<j��<g_�%��j�l#D��i���@���c�?����������K&󾗜��ح�uL�3W#ܡ�q������^I�ɶ��H�HPkGV0��#b�ӆB'���� �b���e�]VS�$ҹ����[V��a��H��t(f�/h���Oz���}s��yW@>�0�����>/]�"J��RˠCh���uĈ�	MV���\���<TR�?����Z�+L��7R=g\a�R�u�(K��x�;�4	�j����SeZ[G���T�}�U��8�T��RPM�P�Z�mo��-ԡ�A-SÅh����A�j2!:���+�"��l=_�!K�������ʱ`�Z'�����X�@ ���u���$yO��$`����7��j�5��&���6��z^�EE
���uZ��e���8k����$���<�X:��$^3q��^lk��Q��gMK��V�S(�;�i|x7^�� ɋՆ:�������2;ٷ�%8<��F�;��E�"�Q��a0��9���^ȃ	��<��������r���q��"�q����>4��ͣ�W���]l���$x�U𽘣Be��\?Φ��nZR�3G����n��%�-�+Nx��X�U�?�!��M��qF]U/���'�}�B�c�>��������~��I+�����}�!_9���T������{�n�;/���
@v����'��xγw�N�ۋ�cY0���p�b7/�������8���ʮ�
mB�^�I����c��C���EC�]��x�垌�w	�p�/Nv~�v�Y<sc�H��$����D7h~?��=NP����}2�V<J���g5,8?���(Pp��?��E�+MТ�Ϙ{�����g�O=���y�@ʱ�`|6HԘ'� �:���%���9�ѕ|�hfSW���1�Q�����PB�T♸ѫis|�׎����W+����}�£�%�lf�È)u��7He�{lL<X+~���:*,�~�yF5C<�Z�ʱ(%~��j��"}V���^Y ��W�7*�jd!ʹ�[ܗ�6��!w��D��<�Rć��;�5���e0����'ߒ���b�s�|'����O]���(���V��@)��'�c�5BwM���Vy=���M�'���i4ϭ�j�{��׵tY���������� ��5�N�:�e�r`���f�ڈ cO&�����~����,>�
��i� �D��*)��̲2c�4&��[i��(�Ƣ�Z�GD"G؅R����|P���]�V�glΏ 1s`�n�GfI���Ѐ�}�c�a��I��Oq���`��+��:(�)F��i�9M;�O��2M�SE���oEs&����T��dT�fŲ������儑u�!JF�5]��t�R�rR������-���o�wY���8j �,�zB��w����+^Ɣ�0��`k#[ˇ@�va4V/xl{`/���m Q�E��y2i���0	� �W���SV7��Θ�l���
��CA�����UKKSg�L��ڳ�2���[�>;O��7N�7�a�js�m���1eG�/����n�a^�����ɖ�ײ�U�ɻ7"	�U�SH�o��,�x^���֛�7Ź/��Ƿ߇��6�,ޱV
�^`Z��}�1;T��|���
+�k���Oh�����~O��;�8����k�j�:_�� F9��`�.�(�b̅�L^R
+q�w&��k�`5;U�^��q�~o�I�Th�/s��a�
�cG��) �B�-q��].�~*�@�&8�#�gb���_�/�������0�U"��S&��/��	����yv���n���Qx"�^i��ܿsD1+I}�D�g�/<��R=�+dz��mȍ���7��s���܁zJ˄�'�F���f�����}W2��	��C�LFf�s�j	~,.k-BE~l2+Vlc��0�ɒ�(��yӦ�)oj�K���&E��˴���6TCLZ	a����.@3�K��9�(�(��_Lȴ��	�3�_f�@�A
������P�^��G쭀�ED��r�~�qi�lA��3�߮�X��W�$��s���a�S�B?\��/��2Y?t�29��H)dK�1�~�Tj�f���@h��J�6J[K/mez^ M�|@��hMs��{�g���,��F'��85���Uwzը��y�������z��"EJ�>-/~*�:�_tE͏GD���E��E����pkkI�~px7����(�)��>� 2h���Bj�⎇g�sҿ�$P��4[� L7l�t[ֲVU�rf�m��Jͼ1��?S)�#l��Θ)7W!����{�Pr~Pm��Ѓ�Ù?�&�S�P���9Se�鷟"ib����6B�Ӯ`�U�zF�9Ӧ�Q++D⑗r���ށ��.N�$?�E�8�	�-���-4�c�kp���B�,�P'���6}M��
}�:���BlO���� �)$Z0l����t���h�K��Pؠ���^xfxآw�|~���BQS�܋�>J����4��xGXS��ъ)Ajr���m���ǥ�e��6�M�fTU���� �I�#i�����*�b�����A���\�j���`�A�>'��0p�A&���S�}�?��wr�45,4�x�ϩ|�x�cB��u���@n.kŎa� l?n2N�����G��\��ָ��������7QZ�B��&h��Ҫ1�Q2R�� �<�L��r�9�俎ZwX���Ƌ�L���������;�~�`ج;(:�P�»�.S���+��;�� ��X�x#�nqg���R�MS�!�|+�Qha1�D��d���D� ����~u��n��W�`?g'��?긪l�	�x>iC��}�e���˓q��:}�$�FV�Y��ЀWۗ��(2�P�:W��b��3�%?Y�n��N=�c(�H�]����iʞd��e�9���n��)���x2��zd2�����Mv<�1�a���;��^����f�4䣜�kJǑ�*����0�KRҩ��m�%��f��ex8�����)�g4?���*O��޼"�Ķ<v��eHUxcuL
rۙ\�vZ�Q���%:$x��{��σ��:c���:�n�>9!g=�A7l\���z��h�x�`#k�F.�+����mu%�]5���5/k�4I��X�����)u9�ɴ��P7��7�y>�
^Vs.RgF��0��$1M�D�N-݉;�p ��~
�����&"O~�=�?��%���|�4\���N��Q��M�Hx�s�b�$p% .B`�A�P����Z6���ҥ��%u�
�jCq�����pm�ý�������֮�H��I7I<v��w�7�įS3�_<�+,�3E�q��&�(Kr�q-�rӯJ3��? A{Ѷ2�(��z(.Ϙ�%�F٫뷹X
(H�q>�Ű�M���@������E��Q�s�4åF��D��)���-��=1V���d*��q��@eX/}T��9Fbl9�ak�$C]�VOs�P�O�>�9�*�߿�n����PS��Ĵ�4囯,I�Y0l��/���=����l�K���Zf���3��i���iË�N�̐g.U��s� �u!��;�����R��Czm��OxA2#�^{���BF�e������nI�o��k�-�/��wy�8�6&�;�?<�z�O 5�_��ߛ=i�YJ��.�$xݠpG�tꨠ�1%�?�
09���*IG��Tn.��.'�2��m���J%�$��[A��)혆K�؍��)� �6ȴ{��.l���`>5r%�&��&|�a�xCROƈa�{�*X���(�#�3wT�s�=�"Z|�w�����N��C���'��spΚG�hScP�S5���.��⧧�[g�@��t^���'*������ �Q#à��j�׋/���`i��<��R�ʼ�FaW���emq�ȵ�gO��ɛ,8��i:7�*�#s*�Jߏ���Mb=[�N�q�@���R�����a�̱;�&B]&��!B����Q�A�Ҳ;/%J��5��۫��;��l�	x�υ�Jy���U�L�
�0ү:���[��1����5�1�!®�g |��Z��0AJmB�Mm�������Ss�~�|�֖�џ�\�'M����U��;m;��	p���Z��ª�Ό�"ЙR(s0�a��3�oA�O��t;�����7��#��Yx�K�j��_=P_�drp/D�U��q��%3p���q�h]N�G/�S���f|m��ב��\�������j�@B4��uB"e�Ʀ������(�#�d:"[����X�����{������^=����^ks4(y7%�@o�PU��"���+�L����tF��
����6��&qT_���E�8Д��-��*?��^���IK�+	b�6#F]`_;�})����ˌ�v���:�ȩX�����.��[����,R���3<�ϣ��$x��\>�˪�U=����qM1�~�M��U�p78f �Bp7B�sY���(���KZ6x}�V�?��x����ߪ4��%>�͹��!��VvU�Y�O�B<�#*J>9�^`Y����H,u�v�uϮX���< r�I�*u��[��٩�G�s�@�I�ma����w�L�xA��8�:�l|Ԉ��ZecBp?'J�a-Q>r-�Q��]��	9��C�˃n��>`04�IP���N�\8+���G�xZ����/�gӣ�!��s�O�Q�@��w�P���lln4"~�8`Ko�38ᲞZ/ҡF�����m.7�"�S�<%Z�������x�Ų]�J�M����骅�[Ƿ��?x���8��8�(tK$�Q0z��X����S�\͗��L/E-6?��f�mj%fc��@r�a'a������.��αwd�T����%m�7��� ��6�H��8#Vy�'0���Ɗ��'#�Ӏ�C�	�������K8Hދޅ����3��7z�.�����M}�/�ԛ!�I�"��#b��M)Z�>
z?a�
n'���yD�Fs� �7��8�]_�ؖҮ^����@�5̻��Ǒ�*m���)�q:o���|�m.�<k��q�k��E��ia��3S��e���N1�K��Ks�����§S��/G�3,���&�C4����������a�
o'�����2`�(��vl���-cƕ�<r�ɘ}�~�nJ)���'��TX��v�)K6�~;џu'���F��{&���f�yPJD/^Ch���ו0�U���'�x�O��~�-K&�3�6�;��[{�?OA�M�O󟄬	���|}`�w��l�>g��c� �5����pY�h�qJD�'ϚVK�Ec��-��~>̿����)�Dk㤃�l|(���de�B���tn�?��In��PV�'.0�^�g�b[7��I����5g�.�q}��D)�1_�<𷬬H��n�o�;Ӯ�vdPC��#T����(<���;3�2d�Z�["������_�d���}#�f#�g�@�?�e���]���b���A��G����'/r�֗_�����8������TW�;�IY��*����������j�p&�A��SY`�=�����%��iQ���V��-����N(�_�`	��U�{���{�e�A �b�Hs�ۛN��'g���[�U���[�N�VZq�������� � �:�<�w'Q���b��	c�%P4��>x�cC�Y�D��� $V�W��G�P�0���60�x���㍶J�G'���B���)۩F���l�e�13	�'�O��U�0d.}W����0��܈Y�,�w��}�߫���v̰Ui}�|���(�G�����M+zG� �4�$�#�uQ`M˭�R8��P�Me1�A1��Qq��/�{�@V�[���f�)>?��>��Uh"U�D�BM+�k���+TB���<�SG��e�~���)����p?8�a�{V���7��a-��҉�����$X�S/�ٟ�X������'��|M��;D3����^��m޵���"� �����H�p�Y\
4�d0�� ��֌daD��Ye�x���`��[ynمP9S����8彷�	�Q`�
E�f��ܖ����A��@�紴�b������j�2�jq��w���,-XfH�1
�1��i/	�����i+uP���T�t�#���	ͺ)d���7�V���<$���@�ǐj0�7!����a ���\�J��9W���n�+����.>��b���8�*4�2͖��I�IIpҾ���:`�z���Ԉ��$��%	;/�B� yu�Po�Ύ���[�q2,��ӷЪ��燯�Q��d(��A�Θ�a@I����=�ե�(F�e����0Wo��������Z�m�Qn�����k:�b���Z��@l���o�a{�֡�=��C�Ԭ�y�|V�v�_�V�EN�7h8�\~����d>��O��}��>9i�&h��V)�q�Vt*���r�ޫ��hڥ�x��\]PJ��.b��T�h�\�� ���/�$�'I�2�����Cv!s��[O�3�^�tnm�Kօ(���%�z�)�F�T�J>���	4oEa�JS��3!�.M���ű֘q@���S�Y� �Q�l?U�6�t�>�d<����D�Q�h��E7�w�1�A�fl~�S,T�^��i��v&5&\�:7��:?�o\�Sdd���RT��X�8�6����j١Ӗ.��.\���#%TP�Y���|S�8������e�֡��U��9����Ib�T�� ��p�qS�����y�'��	�C��m��w��c�:�Dh�E70sn�pP��V� �d���ږ*��]�$'#z�gl�OG�Ɖ���x�t�	U�FZ�tP|NX�^�c�dd�~��#vsu��/�I!���7<5h~aK&�b~W�SD���'�kw3B�[R�D���TQ���˾a���څ
�z�P��!�(#�!A��
'���w������Gy�?���c����F'��KK-���h|ݭ17<]����*�D8J8r~&
J�g
��4���렧��({�A�傺iGy�2��/��lȽ�I ���"�u�D[����B��ϑ� ia�0��Ss��F-�;���]���#VM�|��L�g��7촱�e W�2>s���^�ͬ�ޏ����v�A}�L�/���l��;�z��r�u� �$:XQ��U\��3���D3Ӧ�wf�.�*����E�j��������_'*ٱWM���U����|l�`�O�g�4�pAU�)a���&� ��p%NG ��0��:-x�L�I���/���p��H�=��,�����DO��6ڳ��j���$��X����u��]�d8Z��$��#�f���Z�3��1+#-��U�E�֘Q�;�|�@ZҖx?��Qm�i�n�B���P�q���Peq?��q��~���;V�H��|G��Qp���w�c���JNA�OY��>� _,4�>��ܹ��6�_���3\'8bڇ��R��a��ג�WӞR �%�P�-*Ra�U[��`�BJM�S�����c�ry��� A���nc&h��yMz�S����I�}X��KTZ��XM���W ߐc�z�"��âp]�_�k3�Q�&�f���V&jkV�ٹ��Z v����ܓ�J�����������$�<= NߢÀL#�Tؗ].�)��4O�U���5���y��f�yi��c�x�����]�95Ӽ�tb�A�j���Yà�sc0-H�(?�"���.��٪L1H���%G���ָi�L�LN �U�	y�8�F��	BS.�����Q��)��_|x�_iA���6��g�y����uQ���9x� �-YTXv��S�����,�S�,��ߥ�{&_ekڶ���4P�KR�3�v�D�}�%А\e�R�s|�C�S�lE�2��
k)���Ez��Mɕ-�1���*�A��3
�J��Pr�DW!|g�^D��<�9�l�8��� �˞°
VD�u6W�/p��N퓽E��Ȼ<��v��Kj��r�! ���=v_,9�@���e����4F%stp���P���"/�rQlo�&o�2�o\zy�4}_4�ͧ&#!�E��������x6F���+�i+EJ�2�O�Ԙ���b��"���D�Yk#�/�4�w��Y
v�F9o3��w�#`ψ���\���djas$p�p�P�I'�]�K#b �c3G%q �46rx|��_���jPߙ�~ĺ[�;���/�i�]V���澱����mBi���B�/	k�������^Io�>�M_C܃m�붴���\�'?�4Nx|m-c�U{k
WWu�KH����r8�V�T��V������l�J�5��be���.}���RI:�ͮ���O�C��wX��C�W�C��d�,�w q�ʹF��c�A��1��f����.k�ω�k��ϱ����,�AN{>*�Ҙ(?l���w���"w���'�N�궐!/��Z������XT. ����Ch�Z���8Y���b>���#>q�~���11 x�d������Bl���������25�W4�ї�J��=��J<��,~:����hu������ZW��*Ɵ*��؟t��]��Ƶ�!a3�ᗯ�_���#G��h����/*\aUuhzZ�u P�p����%%uO�`k��`K������:vj��%�ɱ��T�03����~�����4�V3V�qf�"L��*�xP�`�R�6��iu�n3�6;IC���9Cٸ(��v�7OWk 7��ɖ����i��
D��A��/��.��W�� �}�%�m�֢��}���p�����R�T��!��D)�r.�Q����DY�0;��Z9GP���=�βq�E�Tgwc"�@�J���o1�q��Ój}VfDr�9rzϊ����G�[��9��s���C��`Z���v�c���)�W#��)C-�t>�(	��޾���myb���d�&�J]V�E��Yh@R�o�3����¿��x��Q�Wb@�P���U�q&M!;�ߗP1��g����p��&J	?^�C�JUFA��	��X�\u���l�0V�M	�V/z��z,n	�����X9ֵR��KrA�N!���[(���?K�U�2	]6���?x��T�me��!���FY�p)#+���;8�nl����i��x�s0~�篌q���uo8��LiGV��Fu_��s� ��a7�Ua-;�l`Ͳ���[<�!Z�fZq��0�b8r��Υ��ԿpZ~��F�ܙ5xF��K��6����X\j�!}��Y�~|��"��u�f�L�R��d�z{ � �S|Ĕ�;y&���w�'W\|��� ���y���©w����R
8�&�H'��F����b<�S�O)e��*�L������{"$^�d�H��[ �o���H���	���O����K��O����$�슣�|8j�����ia�ds����O-n�{��Խm��:!�^� ,�V�:T�0�$c~=�'��B���޵������$� գ$��Y��>\��Y�ߢ�_T�r��j�aw�[J��/XŻ��(�g$pN�06�r��7i��!X�O�Mv۱�@$ik���Rj1�>�rb�� A��<�x�ǂ��L/���:����mĄT-
@|���q�I_�p�
�9D	��V���Z&#&�Y+j�(Lպu뜅dv|z:X��҇�5�i��W�̿�W�8��G4ỏ�ΰYzBD�E�t(b���i~R��r�U��Ȭ-G`�J� �,ߡ�ə|��vX���7>�&4���%O���a������?����7����
8�֬f;�}�$5������"���ᯥ��Ơ�H�R���Lim\.����لz�>����F��c�vD�)���B��p�֕�5��e��S�����c�"�]b-$+��Y^I���0Ib�#��oa>Mb�u:\��PT� L�;��hYH:mKS���x�� ���s���L:IB"�BK�`0.���]ؤ�'p�h
�ƒ/-����_]'bf�����f4}u1Y��y�a�*��EC��2��w�ė�W_/��N�ru<	�7�0�R�����Ӥ�Ik�ƾC+<[���M�۞>�3=y0
�����"�Z)�H��*���9�5���89���7���S[��h�S��h�)�E�죩4�g��M{��e��c9�nF��O۵v~�l��k/������u@��hz�3�� A�Y��J��4���.����x�""`��6f￝��Ta�Vቡy�ظ*��	A1ʎ�bZi�%2�;WI�7f����R���QJ�x�HA2�iO4Y ��� �u��T�,�~�0�y���������W(��Vx�	m̱��hxtQ��,���.4���S��h��ȅ��-R�	��D"1 sC���n&�oBi�>	���e�)nsC�=:���$g�7�){�6��p�Fr2S�q��˟���5��2̩zM�몤؀l�rb�;>?M��3U�O�@����Hv�(aw��}f��1�>�����Y����	2�g�޶M2c-HV	�ca��[�j�6
�F<~�W1�Ө��;8��UhB� �l�+ڜ� Ohn��ш��'���x�>{��`Y*֠�aZ����k�ؠִ|��!���a9�!mq��VM��f��Vф	'E�c�C~I�������<Ԁă���b�	���1I�K*QL����������.�0��}�ztV䈯�:?�k�e���jnP=9�]W�����h�+�*n��`�Ҝ�ȋ���v��?���5/=B/JCImh�@��q	��RE�+#��݃�,�a[�!�m|��-��դ��������z�x��D������w)�7{_'�*8o���27m^x�i���!H$�����d�˫���ͱ~<��d�.�|怶�D;���U�PtDw`��/C�ܲAC�h�2�%�C�:�2~\̋u���GzljyR�-��PR$���O,���]�s���(i� ��}�2=�A~���X��+���Ň2�8��fDs��Ϧ����/��cV��G�!ш�����BBg��GM�bt*JV-s�!��-�I����	ڍ�=�&1�Q}e�O��յWq�0�Z�y�z�T@}?2a��|�n�:a���E�f�U�J��r�+���E�7�d;���
�2ߕ�#�v�w�W�G�O`sa���~�xv}5pƮ���oz?;�D�i=��PI�)ܐ�Z�9�״��[����싡���5N�{�[ 3��
�'ۦf��s�?�nj�Pd��< �Ցh=G8V�'?���0�K�~8b׺w�ٽ�(qOq(���؊���X�)�GQ"�o'/y�	���v�X��Of�� ?���С�w���]x��Lx�k���L��jU��[,Kg�Y�/?0�\�)��<�H"'o�5�,Q �x�A/;�!�������&���� �L��7=w	5�O�� Z��P\���݇��j�s��D3��NꙚۮ���M�ɻ���c�)U�%̇��/��D`�<�^���M1d^�O�&6) �KhSۢ�4���v�'���F��'���"|�Ib�u1�)��`�`?t�5#1��k�5��]���2la�*�h9�0�5l����ќTh���&Xi�ǹ�� w�$��k�Q+��v-�e�?���A���_���tg�v�O}��M��gU0�x*�Bn��Q����=r��\sB�=Eε�B��2�t�A��MDu�|�RW���^D_��r��Ē�z�ͺ�[%�_Տj��M~�Ü�H��r�]�7�V��=Сu�qe��3�����H��o�@��G-��<o=ʹ�u-^J>��G8H+���~� �go�2w"���K{�����q���w	����[3��<��yB��.��)����H�0+�sjΙԂrLp��RF���H��G���>�JEin�9@�uƗ88�<|-���������G�w)wn\�}���ްȉ�ń0�]�� h��m���P�J5��;��ӳ�}GIS�?��ߧڣ��B2�Č��;�ҳef3$�GD"�3CM�������h�o!qk��`��>�Z�) ��KhY�2���h{J�׀/&�����Y�P����Ow�m�9v_��^d�nR��i1�>+�X���1����&�����%��� `��> �Y��
�0���Ϯo�q)k�:�Y��C���	-	�g���kkk��0��<�����ߎ�OR��$�y�v|X�0F��T5C��b)bȹ���n!�KY��+�O#���4�`=��ƯBNIy���7S<۝�����>�8�����	�S�u���Ն��q����?
�E���E9�:ZD��.�Q7�٫�l��da���
Ò��;Z�W��\�.�<;G�,�2x�i�������W+Nwl�#aű����cY#��&N4c'\��b����>����QQ�ű�ƪ�Umw�9��r?@��9�IqN�K��'��Y���O�5�_O��R�Z�yd�N�c`M���p-du��X%p� ���$b(�z��ao�Z��*��n�얈�w1M�����^�0� }�'|�wʸ��5sh��t��V�$�<4��%(`G�]��> qvќ[69%׉x���b�7�2����NB�)j���B���a��9*�i�uQFэ�a�6H�i�/�/G|�R�2H9O#�)�Hː�Fc�A_��3���G�S��<�'�h,j��l�n�~�}�&��7�ҧ�d��#`��[�]9��kc)/b�F�y�m0r�9F�B��M����)}jc5�:֐h<x������M6|>Z\q�5��[���3�X���,���l���)���F�#�69�o<JL���;+�<m�q5T�#u��S�Ơ� 0!*��"�c{�Q�D��Y�`��C���W�,��(D�=��2k$�̫1<_R!g����
@�r��Susbx�kPeѾ^! B]��
����C�"UT���ن�/j~>^��E*t�vK�u%�Ǹy����?�9�vb���[?�0׽��u��{1n��^׭���ʁm�(��gf($�g�jZ�F�}��1l|I��Od�ϧ/_lE�}���1S�5��?�#n�tfX�ր�Z��?���Z��2��H��M�����~qK��4gy�n���E�[D��u���-���l��D_Ão:<�Y��B�}�����I{O��8�ǘL���%JX��0Vi��kl@Yz��K�sM��~�&53l��p\1�DE��3^y1��>�H����{��k�����#��~Š�6D�5A���^	�I�i!߻k����I���[��]���?�ɂ:C��r�\kI�.�iצ���x@�^��<��J�'��wd�-i{n<밻��-��fO或�_�Rʶz�	� ��%��I!�t�L��F%+9�0��1���<��ᔸ�O��Q����p�DPv�ŏ�A����2��1%��w��#�+)��b:�K:˒j�q�K�`�g����܋B=�Kyaxy����֚��i�c�a&�����M���Tf�� ੺
�K�y}��.�ڒ��+��wxR65�u.V���'$�J������Z#9���m��QJ�Ko�fZj]g�Ǐh�T�fU6\ �>��s!���!QH�p�)a�	���+G���b�� d��yL'�wf�l�3տ�ȓ�e1I`����&�S��~�2�8?{J8׃����^6A㉝R�W�Y;��!�1�F��43�L�����|w�銭,�%ڻ|Y�@���wH4R[m� �o��_�\Gp�ʆ���b
���ݨ�kY���c�g_�o.jD��ez�H/C#C�(
� W0����L#��j��U����F�k��Z%mș.�ª'���IN��+��A<�ѩb�fbLL��/R�kBrU��E??f�������6�<�
�C����rY�l>��?5[Y�=���j>�U�����2٦������ь�
�Zx�����טS5s�g���+�w�5\)�4�B_�#�i9���� s:��Mb5��/�~F����G�G�Ǖ�5��OI��Y����D�O�[�g��'��)�6����?܀�;���NT����+�!��,�����a�2�������kW"-�Og��۩ꃄ��&Ͷ�Q�T ���S��{�)Sa���kI�pux�%C?�B�<��.r�&��19��*��g[�0�D<Y��?�Q��V=�󊕩���!�4�N�ۮ,�*^�6S%��ƺu)���!�.K�M��}�b?�Iu8[�?�579���B�N:�#1���U����w���}�{V����29ʮ_ʛ�i-�;�p�砝�� *8 +?_\���'d������+hB������Q���@�|�VT��!����#Uӳ�W"�ɽ��F�O ~G;��!-d�4��U�.;��E�����wp�MAi����{�=of|�;��"l��z��\;Ӡ8���F�_�g�R��i��м8�J��RMu�i���X�?��z6%�G���͂/�,�ۇu�x󋄙�=�����;(b+Ϣ=���6c��%����~tU��`�y��V.ezD�a|�����:�tW��Mg����z2�Bu#Q��t��D��A���"�R�LvW���U��N�e���(^ST�]���k��Y" gf���4����I���k<���3N@�jǭ^���]��u���!Յ��¢7�1˫j�0!%lv����������֤O��g�,F�l0'��n��U�k�M1#���RW¶���˄"+��d�s��|� ,�;��s�Ŷ81ˀ�����!Wc�v��9�=l�H����B(B<�+ّ.��p7��K�Cc��q�f�"ט�]yeI� �r�����M�DT_6��c�TB<9���Q�M���Cvm1�����V��d�:���<,Ҕ�os.��u���x���� 4�3h�~)�0���`Bg�ye��N�V�©萋/E�$#jU�����K �v��u����=2��j%���`�� +�g|����"�Ck�%C8T;��.�U���1����3���w(�>:=�f�f�UH0#B���I�q���SDR��.�{E7�:Gp�/p3��iVi�D&���3��
������#J;Ԣ6H(�|oZ!����˳+�ؿ�/vK*P�d�@}p[�~y�_~
;���p� 5�Z�`�Ikt�!�s(�]��f՜Ǿ��?�ߏ�-������	�祓�Fy����bڕ��:F���n�'��n�t._��hQ\�V�e�*���;)�y�ƞ���6R9YRʯ��I�i��� �D<��!�t��a����B�I�J��7J{f��<t֏����yĲma}C��6���C�^�`,��}��%��p�;��7���7;-�aM�,[`��,����b�����e׻��������
�<UsN��s����7ڍ���Ыƛ�bz��FK�ؠ����X�q�XE���=�4���U<~S�=U����rYr=j�t�j���D׫�c�f�Q�a��u��UpZ2�F��Rp��F)�Vz���zl����Q䂋Uj��O�Q*c�+c6��<V�;1��\�f'Kowi����8�o�|^m�5�Z�W�� +<����mMrM| ���,9@o��rI�i<kӽW!����6^\��Qφ!|X��#�8�N#���0ߟ:��wS��Q��y}_��d��F���-T#��/�|0�n����e��q_J��̸�n��"��F	3��T�'71�3D����Mz�7ұ�c#x�;F6�>$z~h��W�O�])�D�TAG�w����l�����Fu8M���1}�cyQ�e���>�5;G����Q%�������o#��G�f|��n��q
m�#/b����x:��:S	m�|�Yq<i,���u��{C#�5�o���=�d��
�
�+��>D�!b��$"��pO�O����V@����P�36�������n�\��|�O����*�%���Q�K���c�5|�>Tj ��_����2-9�d�T�)*�>7�I�r�y��t����-���|o?�0w��(�ʎ�1 p�l)�P�M�Z�{�N��Nv8��@��?4��MT�O]��:���*`
�ku�;���S�iŖ�h��uT"��\a���[�n���ӭ��.M��*���I�}��$�#غ���\/��mm�GGS}����O�8@��+�5�A�� �q!�Z���jԸ��E���������Jen��s�b�"��OP�m�����.N�䢅=���=��HT����t��i����ձ=54�S�P��m�������E���������m^�%��\�Ɩ�>���S��g	�����'ύ��T �m$N���$ؼMq��_�j��y�I)0���uv.��.ݹb���z�wB�Hm�&��LYz��/ ��a��5.F��h|���ĆX���0
�9�z�bS�0�{��������'&���z�Kļv�~ȱ����@�-���v�QP��Ӟy[��A�^;����}��-��K��%E��U��^���io@޹�` :,�E�NT��(�t�(�r����W�p�S�=3� 9+�^+�;�RGJ��3�Z-��X�V�P��-�P�6���/�V����sV+�ݐ�DR����Cxs��� ��T�Q�����>7bz��� *�%F�myfqrGU��_�t����X54�A����2z�aU���$�6y_��7�K�Ѕ�����mz�7��������vO@�E�{	yR�z��=��A�@�6���~��'����O$f9�e!L���:�bRy���NV>Xܑ�@�*��)���D��o����8�jhb�$s1���vo ?,r�g������\�����J�o�W��I0�q��,X��K5�l�5]&�r�)�$t2�T���B��㞎�C0��� A��}�An�T���S�K'Mw��,\鶏�N絣4;��nq�?AOԈ�ąe|,4,�
�o\��#�6A�ӆ�_�P�+(��9x�&�'d�9��¸���?��ެc�'���qؚ'�7��
㔥<Qr �K�ٙ�]Xc�32i�_���끧Ym��kYg�x�]�v���5�z# �R
�u��#9<O{���sOuCD���
�^�`��j��_gBT8d�m�r�4H2�� ?�^��F0�E3C?�)��Q���.�T֥	��a���'Z��!)�����yl(�
/J�D�8�K!�X��g�	�ˈQ�Q��%Dxd��
"ܱ��#��칁M�Z�	�-�LhLL���\΄�n_�,�*;봢����b�_So��.��)�⊩e�:x�ǽ����s�~�>�{��Z輀Q@�p��R�uf�	lb�;ϟ8���[��������ќ7��p,��I�⊗��//wk�'����w�Q��*����@�F �:��$ ���6I�Y_��&u��8�-�{��jl���iU!�3>x�?'�v��δ��?`��^�0�QF�zu�0J��3̎$_����;���\zk�՘�!-F�[D����$2��h��.��0g�.������Σgޕ����B���ݤ^��`$�N�S���N�M�o�7�V��c�𜌪���Пn�ڳ��h.¾����ʿ��*�`��q��TK�3���Њ��dx��z�Z>it�b��8�����̩��l�;�����j��Ŋ�U��Se�"�L��Ui�����QLM���Xi�\T��t�`$ts[����9�s]��ڏq¢��X?fo���VPe�n�3a��Z@w�r�5�&��U�y�����킍���8r���j��=��g�y��P�T���Tn�"�"%��_"W�����z��<����o�;S#�1��3�ڼ|MH/eӵ��yu�F
[9
��Wj{�lO�|�;mg����+��#��0�j�$�0^MjD˯us�i$��K�H�6Mc�N���4x�豬L��Խ7����e񾡭�%:�o�Hx7ы�^k���;�a��r�1.�jg�.�3����ZnenR>6(���+n�ζ�>(���G�RK䥁���Z���=�ѐ翷�������� �;w��>���}����(K����>�sܵ�c�;�R�.�����/�S���}�����9�b��z_K��XL�S�^���]P��V`��4�>G�Χ��h�~3�K�����^^���ϥ?��F�gy�}�r��8��������k�b��/��p�ȍ$�`�M�� j|���$����]Yf�%IE����t�ƫ�:)���7���'&P|D~�����m�)�(q��Y2dǖx�21�Ka@we=m �P�F��Z�3wuV��I�al-agoլ>�Ѻ�kf�z{M&Cc�D������u��IY�B�E��w���{�\r�z���M؈;&��{��| �g�Ϧ{ya_�s>��-�ܾ֢2p���P���v��]k��a�������-�m�{�3��D\N�g�ݏ��$\���=vt_�D�!�C0II��g>1�'�Z��u����b�T���k�y�(މcD��k3al�3IW�݇*#P�}�A]@�?9�~�{�y�v���#P�!<jƔ@���}�1�4#�h�|6�7�~v	>��"�{�ͣS�x%M��8�+�ԓL�0����=c ��ql0X�3���z{F�Ɇ�8,?���ɨ���a3L溳wK\��S���&J�*���.%Ɩ�/�M�YC�7���ss8��7'�O�i9"T��b;���c����(vY{-5�cCӦI���o�xj���$m&j8���1�����&�8Rdi�R�N����g	y�0K)2MWZ�J��W.s���x�޲vu<+��&��X=���r�3SM��҇�x�J���B��vQO_ç`?��^��	�4�@0�NhɁ��e,�ჀR�zO���w~0GWwh6�)���vJ�"�TY��2������s@�X�e���� �W�D�%7�M��_�D�$��#E�� _c�&��7� �[/����S*���A���� ��O �8��1����p�/uf�x]YF��!��lAWn��~��[KT�8�#��J��'Y�Z���YAm�Dfޫ���­#jWQ��_runO�����-f� DՐ~�=	��C��O�Mݮ������<nM�[ɬCy����|*:��t���cޱn^�U�"՞���M4��r�=m��L���}�%_����_�71�u�?ӑ@�P6L��p�f�VIH������!e��8���<� �C6�ӗ���2�GV���m]�g�^��f�L�q�20�HZ���ܔ
�!Pd~{�(Rę?�l��|8��|�a�r
#S锼>�`�ͩo���=���F+�d�;�.��÷N@ "�����Ǒ�?j�#?�7��8�a�.,�W-�K��.*Ix�7E��8	�'����x���:Rܱ��]�i` �4�h�ʩv�ɲ�d�#> ۖ�YϹe��������nr
 %�c������C�O�%��|�{�l8,���O�1�0ݰ(��4�q��:RL�̒,�
�m"�V���h�Hr��ݖX���HTXDW�@���R���,Z�����n>�2���N$�y�q�zPWtitq�"H�y*8���)��i���>HYj��3�����upt�Ǹi8����L�NB�R�-��X����y���[:�1�+�%�Kǳ���Oe���J�@
;V �IؓRO �t��3��X��:�Ԓ�Zm�K6���&%܇��`�{�T{��n,D�4J�X.���#�/Ƙ��b�w��t/�IȭD�y�݋�-ձ�sI7"[rό
���̪h�����Oj �@:�#��-�5�GJ\o�k��P&i�A:Q����ǔ��&"przGN��B�Ş��4�H��rW�����j�P����bw��4�g����)�5�X��D6�^;h̪���4ky�h���J�c�� w5A������h��d�X�_H�O���ͷH%��;T<!���OD=���]a[,�[Qgù�|�R�ݲ������t��`��hҷI��{��[D �����n��1�l$�����v��E�3W��*�:#�`�����#A|�mk��������dO#칚���(ڌ��+��ٚ���?S�f+%�J-���Ǌ-��-E�5�__eEy.KL�3c���@������e��6��cGќ�
���h�hk��C}zO~�ݿݢ�O�mo�F*k|�2E�J0�o���1�����>��'�������K�e�9�1����=R�
V�.4�<�-�\������y�c�x�����#Ŭy9V����r� ��0�$A�n�/��2�QdX/�q�\0��������>�ཎ�_���c}q���Ԭ�d�ҡ��6�!̍��*��Jf ��c�ߪ������;߻�}�+"w�x�Eǣh��W�R{S5�.�&T��H��~e�/��K�V~�8=-O�������s��44�]ٮ��q��� .��������O%��ČT�=�Y�,h�&�r\��H���H������C=9u�5�Q팾�-\�2�p�⩿|wI/{~�	ˠe�9HU�j�	ϗ�2��Th�z�K����[���8xw������&E�9�ag`u�G�![['i
��hqy۔�e�����;qyf@�ت����2w7�g�ٶ>S��ݻO��5�+}�����[4���E��T�F.��D���Rt	$�&=\�F�H-I�hjo�x�6��$���L
���J�9I3
�^xhgn%!��X��X���\{m�����Yڝ��Y�����čg�~���	�b7����h������ָ�Uf�UN\A"��&���jE�l9��;&+�w�'��+����#e=n�r���DvU�g9��%�X��(��qժ����#\�j���`�+/�H-��HH���"�&��}�d�T�V�(��k���J�0)�>�O�+�-%�qL2Q��Z��zc+�L�^����x����㗀$�("�՞��q�ZP�L���t���v?�z�d�1�4B���EUn\���v�X���r�$��]�"(����l2�,�W���`�K�d�ܽ���-�U*��l`� "ח���A{��LISo��*����P�<�㡉���߀���:��n��6/DNw�`D-��*�����`�ث�c)�H��S���R63}�����������Q
�<��+I�K�G9��uC����g�5�}!%��$���{E�Ȫބ�;��D�,%��Rcz֤�4����������1�kBlHԋQY%vޞ*a�zE�v�V�ġP=��D.��iz��}�,�d�U��^j�'u���j1�]��m� m���![�(<�> _u�ۂC$���2��O�Ҍp�#N־��j��v�ן��h�+�g*���,/u���|NQ������V�X��.������ȉn"��U�{�Jx06=�P׌<�c��H� v��&Wer����!!��?+����/���q�����Q�L_0���6j������F�wFbh�X�)|͜��!�$tNA�m+�G���Aݷ�Oc�����N(�%e��b1(Ќ�$�q�)d�+?�� ��)�KlRO�+:RӪk�q>�|��Od���l�"\K ���� @D�q<'x����c� ���97�
��&6{n��[c�1]�� �r�q.��E�Ǿz.���5g��ǉ*����
� ����cl~�{{��/bݑN�� �fd�%�ϛ/_S����ms/��?}i�xa��*/z��˭��Ȝ?;nX���}�%�Y�h+)�pBrY�|�F$J����(�i(��#-VZ:X�JZF`j�	����s�
ys��m	x�r�]���|ޞR�Ҩ]�'��* �85�"h�"��U�O,Z�Z���(���NbV�4�{P��O}Y�>i�}W�y��M�q�T��eö�ļ�g���T(�{��*$��9gn�C�2Ɋ��D�Om�T��K�W��Z*���#]�MY5�@ؑ�4��K��ڂ��e2���,����� T`ǈ8�*��l��_��(�9\�EY[�,UZo7To�- !�}�8�!�u{2:1>�H������	�����k��!1ӽs�.���w7��Ŏ�6�%��"��x_����8������$R�2��\s�޶�h�Ҵ�Ќ��,�/�Q����,3v��/w�����h���qj&��f{�8����[4Zwq�.;cv�1�9��m2k�B���l�&{� �}��Km�bQ�#���q�ת�8��Yb� 2	:��Kr�1Ңy��Q2�"&ޓ���5��D�?k�`��QF}��ѻ��
�b����r���CM!�1$��f�W(!�[�HhXuX;��>	aB��~�8��zǯ 
�o�� ͫ�OA�LV
*�~@B_���G�$`m�Q�5��6��B1إ��\���Df���(C��1��㜙��p��B�#-�X�p����WV\���O����8����k��jD}H����/޾q���忎� ��r�f�0K���g�}u����n�4Th��>Wc�*T�𬎜g��4�Bx'^�=�~w}��AU�P�eg�������;��_�I�?U\	��F7����+L�����*g�9�pu}D?��c�O���	WJ�-+غ���܃�ʄ���/ڥ���䵍��;,��)����f��}Zv.r�[��דl��&(,BW'`�~k�z)S$%�͉}�u��"�w֑��}E�r��*�[�P7�Ј3�-�%��㳡D�(׌m�����"�_��Qg�偙�e/�V��܆#����!	��a+�zD�P�V4!��;�G�D]Ay�dބ�U��z�^+Ɠ���u�˄ů�Ve�{䖋�NG�>7*�f��@<"	�nnR����|d^�a��Aޕs�"���,yR��g�����5a��_On0S���B7�w�Q�-C}*
��@ޓ�4�Y"�@�\�?��$��;1�5���)#/
�a=pʶ�1[���@*á��z�Kv��/]�%�RmRJ8����!�ӡ��'P
h�P�c���?_��}��hø�7`6~������J���x�\�m�<����N�w���t��JK�d.[�Z(�6�Z$�����SC083�F��>A�4R+Q7�q�ӿL9���b�������ȅﶣԗ����C�@~[/�ӄ�2軗�E��?���+� �bg��3N*�L��Q)\�Z�x���I���L���9�0��s�݇}�d9J-�D�W��m?�W�`�M�<?�,|�ˠ���F?��_�V��k-L�)f��?xE���d�NN��� @�o��l?�vj��~�bKQ�i��=����Ƈ���&���T�"r�(F��J�����P��B�{�ϡ�N�^N0���O1���}��(���;�%�-�	}�=�����j�pA�3Zk���[�W�Us�x�j�S�@�.�����'�:a��$�w±�S��H�yO�r����sdY��Q!c�韋iQ����]2	�l �$?����z_����VA$^f\�I��G��P ���S<�xH��|��E���=���G��T����(�r��C���dBsbB�t(��=VL҄u��R����{D����J��CzA�R�rJD��
X9Y-���4 �P( Y��TF� �zg��ڒ��h�0j�yEK{o��dp������u>a��;�2=�c:�m�����h�fM4)6!`s�g��j&ì1���|��b�]If
��#�e���i���E�wA޺{��WbI�+�l؂[E��r�7���k���>�98%�E��)��~I,	���J�JHS���&����-빁�?PJ8;
;0�t���sX�(z���{�A��@����&^Njh�/�/�E�y�����ԕ��[��K
���m ��֗8��*B���௩�����+|'(�[Ε��9����gwҫM.��1��
����YP�0<�fʰ]U�������v0U���Ȋ��`�u�tү�3�0���wO�җf|�?!���\;��˜(t��WRۓt4�>�jk�cJ��rn��%�c.ُk�0����S4 ��kc�ה�����B�U�j�ղ��ú7fM~v`�5�/�IjOU �0v?�C`�4��0�cw��:8�@=e#�Sج��q�	�c��Z�{��.��Z��}���<Q�gX�����ֱ�"�<5��s�Y7)S�$��P#�����A���MG��F�v��Qם�v��I�}u���hS01�y,���3r�x+��np��?��4�Tq��,����̽���do-�%�^�H�*t�� _�E�#L���5c�t� orځ;�p��k4Y��V��guDn���JCӨ��H)�er[`�մ( ßB�[G�a�D���6 ��v:>����:e�D�%b�β��/�]mV�+��S&��z���w
4��ˇ�#��8	ˇ~(n�̄w\���X?ɵ�d�H��pD��]a�8Z�q�O,�Գ��I.�Ź�7��!�Ղ��i@�<�å�U���7-�b��AU�1��>!�������K"EC{��>�?F���@�Q��:�>���M���}�] �9yό��^%-{�[up�rDwn�L3t�t������^��V�k \R,w"E����A�/��<�g��5U�����c�Eb���Ȕ�Yt��{��{�Ir�g9�|Ƴ�vy4%�7��`��!��Ϭ��"��m�/���t������`K�sR���a20O*���n��O>o#W%��B���A��Op�.�Y�\L���A����3�f��PA������u�#K
@X��M%5"V)2�,�`�N��|R׻�$'U�p�c��p��K��\lb�O����M"���C�F�گ�ٶ�Ge1��Y4��\�A�aT~�d�IL9���������p���\8�%�?7���Z���L~��&.�3����+��ö�	�U�j��xh(�d����r�m:�/��2�ԛ���!�Y�� #��a4����u�,�s��[��"ٝ4���y���Y��_(^��J�Ц����Sר%#}AMP^m�ITd��>��ů�M��_7>�.�ua�8c�N�é�� �y�a��r�]�A�����\�o)Dy��]�c����z���@K�MF�5��!򟇳�g-h��sQ�7�v��	<}foX�!��g}���!߁/!��&�'*���m:>m��c��_kZ��84�,Rl��ш.��U��6�ɻ-L���:�7�<Qȫ3��B���
Y�@�K����o��#|կ�V��>I(w������5aa>�>������{���:�ux�eGXrӰ�N�/�����5��v��5S�W9Y|-T8�Y��TJ
�@�k�:�G�%�c@�[~K<w�.�h͇U"$=,L)�t�����d�O�?��T�"Q�ɳ��pmg,O~S�g�Qp��T��h,w��̶
e��������h�gc*�aAV�ݙܐ,�&��M�m=�־%tn��ڳ��s��]��<yD��9z��5�T������n�*]s�dL!�_\m�6��oq�	��L"��B�zP����u�r�?�~M�K;zP�͗T-*�&O����������+���	����Ut����X�!�Q��Zq�5��۶��-���	�)�/��?�	���60��m�?������Ɇ`��9͊(>��pkF�XkVU���ca0��k��E�!vg��i+ �����"P-��-N�v#�Dq�����9���v�t}��(z�7��U�y?�(qbj��L�j+���ʸN�����I2:���T�p8J��w-�(ҍ_S�d_��6�8�[��0ѵ���zH� �я���Յ���C��a%����{<���܊Fy��Sv���=u��v$b{=���y��Y����3z������L��?�9o~�EM�c����VX��Y�g�`䜔�X�@��j�!/�6c5�O���՛¾|]��\���&h����$���9�ƕGts�aG��'��p�XV�t|.��#����\�~߮�;�q�����+./�>�e����
FLa��Y�����Z'7Dہ���d�`J��#�3�D�j9���h:б�E-s�V�A�ɽsZ~WӉ�:�ЬW0&b����U�^�,/J  ��Z�t����X��ocӟU.������7P�Nly�Aa�q�~��Hczx�V��i�#bH�U*y�T�r���B�P�/UȎ��,e`#;T�Ȭ��3�Ce�4��ꙟ gV��U ��*@�)xq�$ׇR��2�?N.�CCM	��|u��A�^	ά�xsn;��u�ڦۓg�ɣ�=�e�Y���'cp�=��`���1�"�Z��YV;�=��淥�x����Ƶ�vvDm-n��G!i?�l�;��>���Qh9�s@�t�
���$������q�	��f?.���a��ϛ��ۉ;��E�8O���X���Mo~��;59 [d��;�Jȣ����E�Ie���{�!�	�䒘���s��� �.���<���2-���,@¤Hv��kS��F�V>*^]=$9�x֔�X^����qm�_l{����b��q�L&r��u�~�g�~,�\��J����&��O^�k�v/Q��OC=��D ��RD��Ҏh�=��%���# �u_J-�a]��]���l�-J-W(�g�ɚ�3��O�,7!�e�+>r��)�ƒ�yGA�D�%�g=6�aj��L/������M�nx4-�����N�!��[M ����F��K��/���
����#�iѫG3T��s��f�J`�����-ӯ�}�.t��T�MG1g$���6���M㤻�LѧX���Y�l���f�nK��r���ρ���A�;�v�	���/�:l�|�yR� �h���Ⱦ�8c��i[PH����c��p�q�%�k�ݓB���T:�ǣ�u�[��
��Y[�l�#���}��H:�����d�4w+�Bv&�a��Zb��[Z��?ɛ���]�L�=��6�T��1V2�_K�y��?��c,�ؘfF�넆�c��-w�y~��E�Q	SS��?���?��t(K�i��pߎWJ/�Qk�'�8��)Ֆ�;�dR S[�;� ȯ�GnKa}�
U��}Y�3�y��XhC�N�!X������G�)��.�w
w����)��VQQ�<3�
���P��b��3Y�n��r��/Y �O�+�)&��NS�ՙyDh�V+�%��E��l�K�-�b����$��ME"�$���q&��1;�s?͠r�Y��_���L�\w�9��|����[��-T
=p-���[���țX�" 9j��l������02a�#Z�r�W��|'_����l��~J �,���R5W��1z������e���j?h��µV3j�+ �_YL�����d�X�.��|Dp�%-�P�p�&�t��yoY����UucĲTb�MO������fq?��*�?�m|�s�/Hk4��E�aNT֞Z�����B>�0�A=C؉{�#s|��P=�˴��!���z�Emٗ�;#MSRM�Ʌ�F%�.�� ���)zS��+���{��3��@��a�!�.9UU[0�ΎV��P�X?�]ؽX�R���.����gȝ�릚N�����Ҿ�9������S:Y����g�;��Oc��~�%E��~ױL ;/z�&ڃ"?�j8��_�B*>��;��g�!� >Kk����oP�tD���������
�ƀ�C�&�U�Y�`x��'�N,F�pa�4]��4��s�NӋi-@a�A���Ԡ��P����ݴ0�+<��cw���^m� nM��Y��=`���z��p�f���J(SoX-e�EU
��3�߀:L�W�1��{曦��h��V�"��" @ī�e��"�<�B��	a����F�fWnV(ub��XH#���*�����W�[����|l"��v�/��|l8r��CͪW�
I����/���b4�sD,Ȭ@��P��z����3/�� ]e]��s%i�Pu�ω#ШD`�<PÂ��J��)�!���)�e���g��4N��g���Z�]��o��f���T&}��m�y^T��A1�ͼa�]�f�zY�" ���>�;��J�:��o�FV�)����wCe��
C�|�X;7�j<��|�Lx�p�hgwEF\}]W��q�j�4���U�E����mi�����'�Xݕii�{H�"�['���7��^�L��!����9�;��c]d�u;�^�z�D��V?��Jx�4v���M�|Z�������l����,z(ԤU�)<+���
�%��,nsB�9�X.3c��x�Hd~���uL�3y�-�ѷ�7�c�JChXo^�SW��c���)྘c�I����qו����=S՘n+1zF�P���N��a�	��%^�����
�YD���L+��)'Z$�Dt���[K��t��X�`�P)<����C
'T�}sE���	�q9�[$UT.GRBH�&{���p	�K��\�xm��5d�R��f$Zf��\ο �s��Ǵ�{r�	�U��N���nO�m�+>1�3��T� �Q���+����X�c�X��<SZ�r��.�0D�Hk쟾O���M!��_��%���V�L4Q�OO�G��FZ�I���1�I-}N���|�n���l�RH�,�Σ2�V�x�	��Ekz��#$N�����u��`�yp�UY�O.�����7?aԶ��-��&l�i�Nva:�/�����?��������i̡Z�;��A�.�pq
�@��<8�z���d���^�lVg�0a�ex;�:����ЦS~d��Mb9h��О�p"�O�ݑ�"���y��9e���
|-��J��D!�O	�~j�$�]�<�'.�[g�Qaf�[OR��5��b��uZ1��y?��8ѝ��?�ϭڀ��Jg�?Mc_]�|k�HU�{J��g�h�U�EZm,t��f1���Q��tL��H�h@�M;��P����|V/?ji-���8�t�w��~+'2���0VqEo:��j�Tx��ݺfM4U��H_p�g�*�V�S|M�e�lo�8^���e��Jf;�D:�#��g�z'�