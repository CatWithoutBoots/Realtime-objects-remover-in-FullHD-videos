��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&r�F���oh���[ynnf���6_�g4P�fm���(�T���|��~��h-V�ܮv�	݅+������p��XX��"�f�{�L��9D��;9
R�.mt}��n/򊋓�;��$ܰ�y�\� p@e�K=q���>�)(�|�SG:y1����p"�b�����=Y��ɡ'hA[�(=4w�#��],{���v���0���0V=���ֿGA"��w2"6��=4g�t��xp�`*��0%�F�b��i�\T��3�!l������������X��Є�-2���9�d1!��e�B��C�Z���fi�;p��(�����;��s�Er��`�s�f��i�����m�C�&�;�R�ڷ�;y����O+*鴂u�e�]����s󍡽� ��k�<�2��$9�IK�q�!�쥠���;��>qLL���(���>��-eް 1o�U`��6�S?���1P^��?�DU��m@3��{Y�F
��dG�3�]���@��y2D���b��ڃI�V���FaA�ܱM���ꅇ�`�Q��8�L�mJ�8��/$����_���D����=�y�yjI��|�vVDe�R���S��ի� ��h,��l��"���s|��M3oޞ[�g.~i�sՄ���D��!L�,ɾa�~8P_:K�A����A�ȭ��i� '��@y��%��՘�d�a}��ב�^D�vp+CC��93����°ȘEvˌ,U�[&aeOM����4�Aa�<3�5?7�Jk�*q���zdR�p�
��7в�j��\�G���FCb����TS^RI��8g�bW~��>�i�����Kq�w�yN*����qR�̒|$���2gT��~f��N�*"KX�z�Vh���%;;"���P"=���Șs>r�����$�i�	Q&��F�.������i�K{���l\��*�2���pE0�|O)�����7&;����(\Q��R�a5Ǒ� ӧ�IQr���]K�)zKN"��F��ĦG+�o�$j�0N\��+��Vv��~�R�+��O;?B���٬�����-oJ�����XX(��}�ѱ A�y�n���!]:i����U�������c~�K�;��Le� �^vL�DB�p�A��Z��M=��T�s�&���j�z՛�%9RPij{�B�M�C�`E�~Π�O���#�v�Bވ)H�37f:;�]Q_#������1F�ѯ�o���qnSb��J��
���W�㕋4�� �' �Y���V��,�^��*��3�n2l�޽Ü�r\��a�8	l�GG��t\ ��i�W�u��ɕn_K����;�)��i2�CaB��R��y\6�'�/�������+Ҋ2Y(�N�t���G�zqK�9i�<؊���m�Aj�Gç�X_�5  7���`����ҁ����p3T��(FV��T�6|���v� �|���c�7�L��(a>m��$�3�1��ߨ%v�a�c'����%O�K���A���wׅ������C� A�m�f�mʌ}
��{g[-�-)��t֦�����-��=<v����fh�Ȋ�{�e�h+-v�3p.��/�a����J
��m�-�	����C����x"�Y8m+���"��Y5gD�Y�J�T�A�sѧs�7��>�X�z먦����+&\��aa�8t��T��)�TJ]	�rX�~x|��c�[ܢ���G7� ��|��'t�	�>]D�]��z�����O��������Hx4�OQm�l���a�@����dH�<����X�=�p}LX a��W���yH��`Ѐ��;�fW\f���3l��EQޑ�N��3��e�O].���t9��K4m�@�d&��k4���t�1uE����WE�e,��,8 λ�1�&����)$頀��w$S|/k����=����C�ˡ�#+<|���rI�5G�#����c2as.���Ѕa�}������w��-�#%Ν�\I<��c�]�Q��^ q��RR�j������(���BH��b+�	�)'5�@�um�a�]t*��S�y��蓠�"	�2�@�1"�E]��hZb�b�[ϔ�\%71@��3$鋯4�?V�,I?"�űF�8�4R�K��LLiq���dI�bo�xËEύ2L{��7��*�t106S&1\���(�OE��XE�����ĝLŜ�o/^�M�\�3 �,���:��\�(�Q.���!��RfO�W��Wҽr	�B.��ndוƇ�z/VdK�1Q��hQv�;
�ִ-	_�d8�����١�Z�9C6Ϩ�##�)����12����њ�
���o�"��|�FڲG�O���=��a8v��Fހ���N���xX�o�����i���JvdJ�5���Գ�.�Zx�hc.�\ ���"�������:f#�l`��l���p�) �+��0��\A����sP�P����W.�$���uy����;Q�qA�<��R�c�s�i���Td������ͭ�:�JDJ^N�3 ���e0=;Ze����'k�v��u��^�\�8j�2�c�ڒ���F��Q0��zc����l�����b�d��xr_28�Q?CC%��bȻ�hM�7�f��9!J6�:�¤�v&�J���w+�F:^�jg�M՜)��_����b�ѝ��n!E���r�\��⥓/�p=�kA]v��qy�����k���|*f4J�1�]�b�f��i���c�"8Mv]�4���k��v�*�ba��yε#��������fŒ�Ѭu��!��wt\�脰������g��¬�8k�4�¤���;4�n��1��4�v[$Σj���h���$�/��rSW�J*�J�.�ڲ�{��|�(��E��!Ƿ�gb�?w�KЛv7�iZ�{����N��:��}��^�;�(R�)^��g;D�Q�'��,/��[�0x�q�|=f1r���=�L�cʮ�6�Y_ϙΟYRPe#ԧ��QlNwC�TY��?j�3����'|X�7�~M�<�D'�U+P�z�!f�����A³���?��tX�8��GZ;��`��m �ܴi�N��u�D���J-9��Dx5����)�WQA3�Q���#�#NB��z�@hH��r�7�]3�f��:�\TIf+�=�Xp�� ���d���s��I�={�}�����8Ȅ��i�ᜓ�AWLQQ�#�ـHRP�I��ײ���o(}Gt��C�^^"2����ھ��~�^ԇ+`�>�0I�?/����/�Y�:v�%_{��6�3�C�,�ϥl�U�����b�������WL��m�8ߙ�f����jb3=���J�
A�ǳKu3x\�H�~D?�Aj�Pr�/�`/���\���ۏc �wז�,+��q��lh꧝��o�j�j��q���+��G�5)�����lFW��z=�ߗ-, e�O9 fב�c��ٮ� 93ۈ�y���Hm�ë�̮�Қ��k3�^Ȩ��t>�C8Ρ_�m�ݨ��l3�Y� ����Uy������ڕѯ���+:��J�k����F9R��o��,��eK��,�$=�I5׈$�
-�䇯�%J���7]�2�����j��^,ik'�� ���c"��%��{U������u%e+���EKi����z4������}|����B��!��1�H/0B'N���xtr�I�ʰ����j�!<���@tC��e0/�к>v���g��pU*��g%DtR����K�������q����{2W�ߔ��]RW�jyx����2�f�����)~�.��$bצ�����^��B+�������6WƆ=�����u�=���{��X$�|���hߑgn�p�gp0�.����+Y!y����4�Թ����07�Ӏ��� �F������륺�/�FpF���e�7���[1H��x�p�b�y�*hu�{-��`��b�l��U�"g�iu>yp�Ds��KrsLa��R���(��·vc
��W��
Z�D
���,Й�	k��F5&y�J4-ͧ���\���<Ub�E�65U��>M�' �ΧnƯV��V"zV3	g�ݿ	�sj�9���j����'��KC�S�a c9/���G��E���Xu�:
��H(��!�q��j�E�%�wYĩ��X�]�-2>^����������ѕŀ�i^���;�*)��ͣ��Eq�$��qt�tH
z�@����s�.�3�qa��*��p��F5/�ѽy_�Q4<���*���m	��T�4�*uxo���L�O$sw/����roq�����Vrw�?%o1|�]{skB�� ���a��qh��y]���ّ�ZB�9lC�OaM,��$�
�(�*G@�~�Η�r[\���Y���n��R��x9�>U�g>����AUM�9\>�.$�K���"����W9+��Wv���hwJ.G;��^���gz��͙ T�����}���3�9���I���yM�_�m$�(�-�j�9��O�l�}e���/`���Jv��Nߵ��=� <�wlZ]�#vP�.�����ԍ/�z��sB�3��n_#%�;�ui΁&}*�kO��}ɣ��ńڬ{����k%!sE����p�i�K1?(J�t��!6@2 ���9%b��1E��&%Bi4A����Ƨ ���Cc�;��I��u68�O��4��ʀ��T��2���!�R�{���	����vO���B���SBq���6�Gdɵ��5�~�1(�w�x�����Ѝ��Ǆ1��bۖ1�h ����vz��;S6#����kN|�i"ؤ��<aX]Fr���d����{�z_qi�
�GbV��ݴ��r5�e��iy�?�v6��4�ea�Jqŏ�f����3|!�1�M�e�$a�'��F(��C��^�݀%u���u������b4��?6���S���tD e4|�GqB2j��6�Ħ5��_|����n�wX��Y����k�,˅�ԡ�,�������A��fu�����X���WiV+����a��2׬R;���mIVR��}F<#;�fM U�tu�H���	*�e��(��xh��2�ZzT�W�K+-�hMkG�4C�b6�ڰ<��J簑����l�2͔6��۔g���{��n�O=k/B�`u��X\�	 ���3��]��B��37�<90m��!�X/�ƹp�uLo6b^1}�)Ó�3}�j���)�]Ǡ[���閫��X�.'&��&٦�Cm�T�6�T\��.�v-�rw�J�ɟ�U��.�:���'?j]4����\B}�o�ȌA~K��)��G��n)<��]�w9��JL%b�%�c���#[�[�� V�(���,�����Q��z2���=��_��A�K�#�*�IM���S����K]�����)�ּ�DbQ�F�>��T{A�g��P��\���;�vk��f�
�zf�Ӹ�N�i���ה��9M�*J7̭�$|a-��_%�Y�;=�8G�A�g���/� �F�~}���s����aP��ۑ��b<��:g���H���+Jk�&�0'�*�P��)��tu"���^��	���جO��e�s�x��@����[Ξ=�!��0���Mu1{n�ݺ'B�� 6�JHt�+g�-�:US����X�f���}��Amc��o֕'G��#@�����;��LJ��lN��Z�6�Te��3u%�>9�&�m4&��"���$-���.�<���{��e~����p�&�.�ŧ��n�D)�P�ޘ�dحm��ԍ��_j�}9���N���Q�k�֌�jR�c�n���|H=|b6!"W|8)��W���p�vs���ad!��V�BC�>CL��0���ҹ$�0�.��[�1Ⱥ߳z��g��2����f�c7R�>)�2�L.�|DU+�:�?��5B5�����c�՚��F�F���!B��f����71��+�����U��n`�y�YRVd�V�4V� }�Yw�d9�� �u\��L��˴?1��C2���Nj�*�M�5<Ԙz��_TՉU
�R�#S��H:�DjZD��/1����)'��N1!�8pX��K���GO�Jd㗎C��97l�L8J3G�����?	B\mp�5�1�3	ĵk�u�_��7L}at=���}�jN(�D���s�+Z�t�s�Ī�8Ka'jp��x�11�ȍ�W�8D,F
�qAyF�j������Tz?-=�G�L��WNЪԇ�z���C�������̐5�qR�N��o#;�Ni��Jp���k����ʷ���@���ެy�H^m�54|N�Es�JR7�%B�4��b��F3���n�yK(�\:�����Xњ����C[��l��ȶ�X��M�v��6'K؝oj�D���}�Qr���0�`0�?������ܯ�_t��r�C P����"��ܿr��'|����h����È�X���ky��@�Gm�d���QL�8V�!g�c4���/5�(H��t�5�r�b_�n�������$�&FH��v�	D���ڤ� /o��y8�o Wm�v���OK��K��7;=L�x��Ⱦ�a9��.^5���b�}�<�[59Lý��p�0��{RG���j4�H��k���oˆ0���6��\�Ab��=ΒG��ْ��	�6(���j����#���[��&RZ�U�����WJ�֠!BR=�b���n�/|)�0�&�2l�nP��Pz�7�PN"���D�*�����}����*Vǹ��SsEY����P�F�H�$��v��'Й�����2])��_A�(%\+3
�Ј|�6�mc��.Z�y�/�L��@�Mu��R ��aѥ�P���D�e����M�!�����Oa�!m��o���ߡ���G��\�����Qa�FU6�+����0>���S29�n��a�_�2\ܩ�J)��E<8�כL�#��i��$C�m����f� ��E��u���Đ7�_�O�j���TQ����\?x����瘟^��U���>%�r�{vbH�"�b��t):s@R�[��-L�M
���zV���9�!��@��(�?<�6FJ$e9�"�$��M`-���5Pp�d$����2]]�+�V#��%��UR%he3��'����=F�w��e���"�I<?�]�@�k&%�@̜!���Ȳ�������������мgҤe/�,Vh��8y�%��!��L�;�iד�C�D~�5&]YE�"��[x��EM�r�D[Ͽ%��)�l�Q*����G}���d���#:���u�5�~�fu{�=V"џ"�cZP@&���,L]�P[���6Rr�c�W�0M�ϕ7����A���n�SJ�����B?��#9�R��*2��jQ�I�=�͈�}r4�0��L��A`??�3�z&�K�DP�p86�5TP�A�u�[7����ҌRJ�wty7����IV�$E9����	ֱ�_���wV�G�d�%��o�Ě�ݾ��Åb6����ñ��� %�0�V/�ސ+�=�!R��[�n����Q�����J[\1|�n�����?Ǎ9��qW��<�A��ę!��0�7�IP� ��<uV��4�a�����M�z�]�_	�[���~m��47��~l�m��Ij��r���t|�O�|��C�ώ�!��^���r��nԕ@���'6��i>cJg*�K��,x��m�UE\�FJk��k*(��)WzE���r�Je�_�50>��������LAg�]�@e{PleV����� fix�c� ����+�����c�27���8�Z�ُ+$՘�e��B�;B�Z�3�n�~ޏfr�)=�;t
'/mI>�"�/V��	Vt��7�����	hZ���(Tm��,��&]��'�o�����8�����Zʛ
���MG>KӴ��n���U8�����ȳ��U*��V-��uY��Gn���۪��`�b��:q�l=����{<�s���JQV�a�R)�$9+Y�ncgE�_���4����)�	��/���Ƈf_.{ĩ�w�[�ބ�e�?	�*�fh�1N��K�iJ�b~OA�fk�^��q'�t�Ul��5*��������6]d����3��� �-8@5���$��ܲ<������3�o�o�*�����e�rm{,�H�	�s�n�|����(!�e)e��2��ᘦ�u��i�m��gu^��d��Djb �.T&3n�
�(7�}���T�i$G>�}xKACw��(�K6�(x��M��z�r� �B�K����օ@��4K):����;k�y"J�A,�?�oK��3$�U�l_�Ůˉ�Ƃ��ƹc�4���p\�>�d�XY)�5w\��/�P\��px�W��j�pF%O��k�4�t�8��(���.3��U�����0�N�+�>�t4���ч"�>�A���?<P{O���i���Gr7����BY�H�$��z1��C� �bT�JKE�O�!J��h#�����*\�R^�@7g�Z=��k qLS��Hi���(�Bz���2i�߻�g��.5�`����Se~7����ٖ����`&sr\���wQ����4b�����a����UI���sQW��� S@lE��%1�2���u���X�Mg����sjY(�	�� ��1����1!u�L����5�۸�^�����O���D�T�c�"��I��&���Pr&�M/����VM��"�Ҋj~b�Zxp���7�X�3�˩����`^-��A��%����2����e�ƷK"$��Q����v_`��ͯad1��3�RP�����|M�\������q�y2�v�yc�IJS80V��hR�y(�yU�՗-waa,��6�G�-[�����)�d^!B�����ݺ|,��~_]�0A{�ۑ�$��QW�!L�of��8�}D_JL��A?Rs��}�Ze���P���5�e]\k�5&��ؕ~�Q��y;�lw����B���Tb�r�qk�p
�d*6~�8��e����'H��e��-�z�@�؀�c��teTc���=�&h�,4i��Q5x䝕.�J�2��j>o���5!l�������I�-#�O3&#2{)�(��ܜb�aU
�>�j���*/�I��qX!��N4�j,�w/��-��� �IN��U�qtV�������eZ���'@\a��v��&�^x|Sܩ]��r;I�@MXS>!N02�c�T�T~2�a�G=ePlyf��z�����-���0�-5��8��H�3�Θ0u�I=2�6θ�{L�b"��l�H�d[z�9L���AǌMs�q�{�����u�t\x9�P�ƴ9�_������J��%�P{�}G�u}�����Y���U.�����]t�.�Kè�f P>�\;�˱M������4����Ǔ�צ7�]�ZQ�B�i^�i���+�2�/�H3���.�@7ZQyE�O3kz�?3L^nzi���_��/;���e���P�РSGT�i
k_͍1/�-{�k�0���,'��l�I6��Z��`r&=V�O��/���g���y�FTɔ���Xd'!��i��t���o���:0OZ����=��1�"��~E�f�n�Z�i@h&�նۗ�TAf��0��)sG�q�lJ-I�!��5x�vGm�[�W�BΣ�$NrY�O�D8�x�6�� ���FĦFH3_9��Ez�K�Dh�K�mJ� �	�����I?�y�JZ�կL��2\e��^�]�c8ב^a1�#�+:�>�ΏnF⭖�P�8�ℹ�L���vK�3mĸ�d����a��B^�z���8J��Q�Q{(�x.���SbPa�S�!�]��h,?��1��M�l+��#�/�jzV��<�aBf���>�k�^V��p��&��8�:/����j�ZAE+����S��t�P�~L����y ���j�4M�p�}��SYP�mm��j����E?�t51�A~�}��=�s�j������=���9����"���d,���a��p�&�\�<��ڌ�!Ԛ���}�3� �2���/Z�]b�zY�4V��~j�I�U����f��F��W��V���>����o%ܚ��s|� ;�j,�ڢ4;l`�ɼ"��џ\�"�{�����?�����ف�߁P�C�2Bf���Q��B%ӭ5��f��p��P�Gء���ɪ�Y`#'�gųH��f��q{����X|y�p�X�2
�\&�]\V$E�����Qlt1���>6����=��� Ѻ$�� �cЋ����w�kr��:��E^z�4����C.�ȃw?�9�d���Ll��+�����Y�˾8��D8�&�D�R6�;�jR=�obd�l�e� ���i�Av#�>K���je�4H�ЛT���1t�q�YrKz�!�]�%D�֒C�� ���B:q-<	kw3X�M��]y��QF�Hؚw�I>�ͯX�:x�M�&p��eq>}Y�7�z'Q��>�X����
�AûY�9��li������a^�����=�K[��GQ7��m>��Z+�}BmJg�?kh Wf��,k!����]�KT����Q�9��A��7��@_���hsqؾ�] ���W�P��
����J�����ݯ����U�ѕ��n�Rj򏭀��3�`P��k!��_�yGS�3���_��8̀R��¸4��nX\�QNB��f�E�5:cB��ߝ�T����M�3�b;pNM�aջ�Ź����Y_E1sI�7wS�6�8�r���d���y�
�y�V�>�&�z�Z�	�Ȱ�PH����m}�s�4ڛ��Τ$q������5.N[���y�?��5b��֠�����z3�M��˄��|���TҢ���v9�"8���οǫ=&���X��rK�����#��+i��Y�rI�b(_����h{�r�&�J�Hd̳�]e��x����4��Yvlݯ��C�$i�Do�;CءRD܈����P����d��E�޵閃�L�1���O��B�Z�7IUy������˝-�v;^뛙�z��룋sf)�MIzMC��c��^cwse}n���%|��.��A� ��(�ǒ���+3z8�^����&����F�B��?�"�x��!!�o��dF§�������f-���MG�g�k�+��ˑߟ� 8��z�?�9��S����ί���iU�Q�H��8�X�a����4�#��İ#�ǔ�Z��Sx��g���)��/��tآ}|�5���1��`�yp�&���#UD���[���흋ʺ/�I�0\J~`欥�Q�[�K�2z��Y��䗞J�dɹ��\���. ��0=k�AQW��bF�n�,�44G��dJqt�oKG�	������%� �8�O|���t,�:���\�X.D��M Z�d�q�2
k^4�4���k ��Z���Hzd9�7��"�e,c�!@G*���KvΛ�V������.�E�iJT�I���ȫ��/�շw�	��Ķ͘� ��.�����\�}[e��c�_�0������/�Ú�(޲�߮�Ա�7 �=3���_ߪ��p�f�j}a���-�G��Fx��s�2Ng�jmA+J�m�}Li�F� �I���������ު��|�Bj鎒a�3(�,�-���&��cD��rA�Ү�nt��F��:P]��-�O/�~/Z���!��pe?�L?��1����>�JlO{Oɒ�!UeT��y����H_<:����4�����o�lQ�/�H���Qa\�tu������z��M�����~�Y�4�+���<՝����[�eQ�y�?�����X0���e_*���>Ás�bnM�5������)t��M_;=�F��`��˅�����\�V0Q��z\gւ$�T?p�Bii3�Jep��m��w�����V���4_G�4���m�ڱ�{�>$�g��g1��Y�%�ģ�S�Z }�SwN~�U�i��u(|�Xk#�D8��Ԋ�v�4%�°L�<�`D<<�dsa��l�z�s�F�0�_@&���{��ؤ�8F�c��G���P��<˼�)����=��O����Ǫ��m_[�^�&,=;k���z�J�����F��y�k|�M ���b͇�(��`�s���
�z�ӳL�`n��@�−i��}�W-�a��e��X��H^�U�-M�x��X~C�F��;��r�˺ϼj����l� Xm�����J�GGa?W&-����:�c�@������d�ߟ�)���D>�G66x� ��H���1(p)Ar�R��7�iMz"\ϼ�(�k�J6T��G�C�^_+D2�y���F����Pf�x�� �q��׷L�i�eΏ_��>vE���Z/�[e��M��}�Eΐ5b��t��N�$'�6�����0����o�RVQ��#I�l�<ʯ�xsP|�f�B&�.*�TF��ՑeA���k��^�KqЦ.�O��`s�Ƙ�G��_x����t�|��C6M��&��)���⥽�&@�KP�B�~�%'�n۸졩�|��a��k�� ��x��o֓�:E��~;��g��%��X�Rxl�<~L��.�?B
�k��>�l�6`w�;]�HA���q�G�vp'D��Ś6�5c�����k���"}�z|�ul��XD�{)ת>�p1M�	_�yTQ���<�������pwm�
�f�F�6���g����e���Fm���=�M�n47RV�@�5y�)�	�9��Z{���ޛp�q0U��Si2�3����Hړ�{N�k��麺�|*ut����P�i�ȥ��<\߆�(��>M{�s�V��<O�}ǥ�_J���c:�͸-�=��
훸Q���+ڹx�E˰D�A����*sl/c�v��Fٔ�J�I��yI5p%y{�Tϣb�ӌ����"|��k�C�9��3'��� ��-/��Yt���,������4�Nu�1���2��T���Nf���?�a��Xm�0�S�4��,�5R瘩��A��կ�j�'���&�O� r����W��z�~-8淑z�>Ҙ�v�t� �B���Dћ�b)�0C?R.]���$���b�԰�%f����2Jl�o���aj�KgG6͆�=1�3��k�Wla��P�T�鴂�`	�W ��Gv(Ug��\�O����.X��R��JQj��Ȇ�8��T�m|��S9+��tF�CJwR�[�	ʹ���bF)�l<�#5C�+�^��x��C(.L5�2KÄ�r�CqS��qԇ/a�Ƨ@�\	�*v[��6v���x�T���w�h�F�Ӝ���!�xg�~%�6���3;iFN't�gΏ��0�ٹfT�iY�
u�����KP�S}WZ��U�/-���b���ލ���j�X�{U���C��=��!]��:h_�І�bV1�0=yK�F�+/�o���#�M�d �`��+x,�5�w�?����������"g���.hJ�9��W����⭦م��)�%='�{irR��eD"bw#�����W������=G��-���;�)�p��*��i��w�{S���:�_s¸�y�r��!թ9��F�``c�9���x~�T�"�r0��x��p�-L;�0!���b�Gs�`��]�ë��:b7|����0��l9:BW�	��J���;��,x�*{�A:������8`6���	�N1��ua�>�����R��[k:z>U��H��i����*�86����h�3����^�.�o��6���e� 4��)��@q�	������<B9䀡�%�Go�+wA�!wǟ�M�y\K]�^�Q-�jm��Kا�4M�*qK��z��^M6�@P4oi�s킗�R��w��)UpY�Î�
 B���z��8���T+�s>Q����S�b𩀚��cs_���cn;3����bOn��B7�5�����OiR��Y'd0^��M�G��$c�۫["�8⩫XVx}f�������f�w%�}\��|؟3�pq��2��*��i��C<��:�T'���i���a�u2�ZY����"B4�L}����4-~����z$��oA속M�*蜦Tyђ��za�pn��Mx�\ ���ؔ5ּ���³%���K��=)����ly�4�.垖'f�e��{�lKo���q&��G~��#hEo�OmM�S,)w�P�_D�B��ᙁJp�o����
t��{�Tu��p�F����׊�6�S���Ҹ���}a=q)�r�)�/mb�OlH����$��Q�%Ea�5r�H��~G9�b$x��g�KjHPzi�˻��7��	���2U���Qd�1T;^�+�F�	��8�2(�+7��Q���LE�aY��V J�ʡVĕ_�� ���ȓ�����(��ȍ�h���X�PE܀�gC̉���5�<���Ó�,fy˫��zKV�y���
��2It����u")�v�Q�iT�#zu|=�$�@LQ�=���2C�%Wgd�#,�ME��)�2S"g�,D���hI�������2%�
��q�ܿSM*�q��@_2�����˒��S��y���;k�}X��b��D��=L�޾H�����}`�y����VT�"� �C�P�w`Mh������Il�?�Y�F<��^���V#�B$����`��e�hgg��\��0�M��~��D���]p�@��:=��S?3O�_'�z�E�ؚ�~���4W~fL�{hE84X�P�Z�c\��IΣ'�7�"tr���q��l4zms(F���TX��g@{��o`���F�4&w�$��R2��&F���ۍ���S��.z�j�ti��A�����C/z��u`�'>a��(�v+��沗3J����A�u5�v�+H�6B9��P�C�ͅVi���,��("�����!�/q����qQK���
�,&m�A�$�r������&,΁��'���>O����F_2�3���o�Ñ0����m⩬�Ͼt�ａg�>�?�W��6���n���9��wy�D}�L�\Մ�6�6a��27�J�[6���3X5YLϟoR�QD�����6Js�9i�ܵd|�ȢYzXyc:n���п��CN+o�<�5���jE�.�<2��d5�y�!̓*��K���$LQ��5��L�&i