��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���<�qO�X�+�`"Y��KkA��3���C�E�B;y��w�/�T?*� �/�7]��3U����%�R�l6�V����G�l�T��2�p��'����2�r�ć�5販��䤋�4���w7����f�+�۞�i*kصZ���a)6[\�@���^��s}�����^��KF��B���a�����ItQ��Z��w��ol_?��1%	"JLH��5F���V[=�S�` yJ(�$�'&[>�:G���?�{G�*X){W�f�[vM��g��(�����S��|��g�W���U����n���$-�����]�;�I��SZ"1
�7��*�[?����e��ݲ���w�*�^u���%Ob�w,
/QW�:gV��[p�\i�ݬ��<����㫠��x��ݓ�z����X���7BhVΑ�wkm�xR���J~��U-��]�'�m����YxD@�q�F�+����tj��=S��6�"��1nKQr�b�t��l��&N�����iC�y�3Q�^'g�@q1�R��k� �#[{=q>9:�Q=h�/�MzGШ��̃�{�]-���_C&��bh����eL�A����?&��n8� uI$[�Ey�ku�ZL�����?5>�x�b� �1���qы0����/W�É�04Ϡ�=n$���c�aO��x !0��>��2������1J�}VA[f�)�"���dzfu�҈��?�u�&}qD:Rmԩ��-����A�u	+��Ñ��  �&����y���^ �Aq�&r�F���ohD޸ayD��r>���f:�w ÷OU�J�Kv�7fN�M��#$2Ep�<Nׂ���/}e�S	�!C
}℧龵qC�>����Ox[�r�"d�],��yi���#ܔS�(�����y@�4<�~�ji9���8T>�=s�x����>EXԬV � ma�|��o�骢�.���h�l��ﲕ΀�-K[F�
ET�t��N��m#�Ί�t�: ����q�I^����Ž�҄����o��� YXnB!ӳT5��MP|4v����i7ه]����5	bHN�/DB�~��$C����c8��Ƞ;�ѫAE�Y��d���]�v��ܮ�F��!���bP�,��E���P�H��Hoe�VI���P�8���V����
M�пTSʸ^�]>  ��=�`1�����U��mY9&�]X����Lfk�e�,��v�59�!T��fB���ti@G���0_����Q%�!��N+�u����K��Kg��rx诸U� �f�A�(��M��L�k4�B^���6q�̓?6�ܒ	)?3�`]L��i�x�e�"0<n����J�<��]>���{^ �
ŊTn9�@h{DTڻ�Pn�4v�
�����M�8��A�'l?+N]��8;"S��iZ&��;�P!�l� ֽ<�HA�X�k����U��2�ջ��6IF�T���8&P�\��Rg�,<���l�V�H�L��tK:�S������z)�,�`�%�?�Ô"��L�S��л�͌_�0v��}�����s,����$�@$}fE.·�Y�����?���A/��>�uc��=ٚ53�*��څv��cW�NaF ����,����AC�!��g;�F� ���'[ ��4���[�t���p���+�
J�]
��U�#����}@�{�@��h[?r���03�YO�{�Ț��Y��]�� W��0:<��Ѭq����Yy���^��ƪ�3�q(�v�м4[2�&T�ƿŔ,�z
G�ձ�����E+�Kv��=D77ϵH�� 0���*@�N83Nƭ������f�?�����B�T�nOR�.6�%Ǿܔ�����-ulN]l0&�Z몊=a�(py��K��P�!����ɕ�:�I����4���	�(��N$� K��*e��eJ?�_Bs����� �4'��>#
���+���,�}��kz�D~D\0��}bۥ����ʡ�p�,